`timescale 1ns/1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date:    13:42:18 03/17/2015 
// Design Name: 
// Module Name:    HCORDIC_complete_testbench 
// Project Name: 
// Target Devices: 
// Tool versions: 
// Description: 
//
// Dependencies: 
//
// Revision: 
// Revision 0.01 - File Created
// Additional Comments: 
//
//////////////////////////////////////////////////////////////////////////////////
module HCORDIC_complete_testbench;

reg [107:0] Instruction;
reg [7:0] InsTagIn;
reg [3:0] Opcode;
reg [31:0] x_processor;
reg [31:0] y_processor;
reg [31:0] z_processor;
reg reset;

reg clk;
wire [103:0] Instruction_out;
wire InstructionAck;
wire OutputReady;

parameter NUM_OF_INSTRUCTION = 100;

reg [7:0] Itagregfile [0:NUM_OF_INSTRUCTION];
reg [31:0] xregfile [0: NUM_OF_INSTRUCTION];
reg [31:0] yregfile [0: NUM_OF_INSTRUCTION];
reg [31:0] zregfile [0: NUM_OF_INSTRUCTION];

HCORDIC_Pipeline_FSL UUT(
    .InstructionPacket(Instruction),
	 .reset(reset),
    .clock(clk),
	 .InstructionPacketOut(Instruction_out),
	 .InstructionAck(InstructionAck),
	 .OutputReady(OutputReady)
    );


integer f,y;
integer i=0;
initial begin 
clk=0;
InsTagIn = 8'h00;
Opcode = 4'h0;
x_processor =32'h00000000;
y_processor =32'h00000000;
z_processor =32'h00000000;
reset = 1'b1;
 
#20 	reset = 1'b0;   
	x_processor= 32'h0;
	y_processor= 32'h0;
	z_processor= 32'h0;
	Opcode = 4'h1;
	InsTagIn = 8'h1;
#20    x_processor= 32'h0;
	y_processor= 32'h3c23d70a;
	z_processor= 32'h3c8efa35;
	Opcode = 4'h2;
	InsTagIn = 8'h2;
#20    x_processor= 32'h40400000;
	y_processor= 32'h3F800000;
	z_processor= 32'h30000000;
	Opcode = 4'h9;
	InsTagIn = 8'h3;
#20    x_processor= 32'h0;
	y_processor= 32'h3cf5c28f;
	z_processor= 32'h3d56774f;
	Opcode = 4'h0;
	InsTagIn = 8'h4;
#20    x_processor= 32'h0;
	y_processor= 32'h3d23d70a;
	z_processor= 32'h3d8efa35;
	Opcode = 4'h1;
	InsTagIn = 8'h5;
#20    x_processor= 32'h0;
	y_processor= 32'h3d4ccccc;
	z_processor= 32'h3db2b8c2;
	Opcode = 4'h2;
	InsTagIn = 8'h6;
#20    x_processor= 32'h0;
	y_processor= 32'h3d75c28f;
	z_processor= 32'h3dd6774f;
	Opcode = 4'h3;
	InsTagIn = 8'h7;
#20    x_processor= 32'h0;
	y_processor= 32'h3d8f5c28;
	z_processor= 32'h3dfa35dc;
	Opcode = 4'h0;
	InsTagIn = 8'h8;
#20    x_processor= 32'h0;
	y_processor= 32'h3da3d70a;
	z_processor= 32'h3e0efa35;
	Opcode = 4'h1;
	InsTagIn = 8'h9;
#20    x_processor= 32'h0;
	y_processor= 32'h3db851eb;
	z_processor= 32'h3e20d97b;
	Opcode = 4'h2;
	InsTagIn = 8'ha;
#20    x_processor= 32'h0;
	y_processor= 32'h3dcccccc;
	z_processor= 32'h3e32b8c2;
	Opcode = 4'h3;
	InsTagIn = 8'hb;
#20    x_processor= 32'h0;
	y_processor= 32'h3de147ae;
	z_processor= 32'h3e449808;
	Opcode = 4'h0;
	InsTagIn = 8'hc;
#20    x_processor= 32'h0;
	y_processor= 32'h3df5c28f;
	z_processor= 32'h3e56774f;
	Opcode = 4'h1;
	InsTagIn = 8'hd;
#20    x_processor= 32'h0;
	y_processor= 32'h3e051eb8;
	z_processor= 32'h3e685696;
	Opcode = 4'h2;
	InsTagIn = 8'he;
#20    x_processor= 32'h0;
	y_processor= 32'h3e0f5c28;
	z_processor= 32'h3e7a35dc;
	Opcode = 4'h3;
	InsTagIn = 8'hf;
#20    x_processor= 32'h0;
	y_processor= 32'h3e199999;
	z_processor= 32'h3e860a91;
	Opcode = 4'h0;
	InsTagIn = 8'h10;
#20    x_processor= 32'h0;
	y_processor= 32'h3e23d70a;
	z_processor= 32'h3e8efa35;
	Opcode = 4'h1;
	InsTagIn = 8'h11;
#20    x_processor= 32'h0;
	y_processor= 32'h3e2e147a;
	z_processor= 32'h3e97e9d8;
	Opcode = 4'h2;
	InsTagIn = 8'h12;
#20    x_processor= 32'h0;
	y_processor= 32'h3e3851eb;
	z_processor= 32'h3ea0d97b;
	Opcode = 4'h3;
	InsTagIn = 8'h13;
#20    x_processor= 32'h0;
	y_processor= 32'h3e428f5c;
	z_processor= 32'h3ea9c91f;
	Opcode = 4'h0;
	InsTagIn = 8'h14;
#20    x_processor= 32'h0;
	y_processor= 32'h3e4ccccc;
	z_processor= 32'h3eb2b8c2;
	Opcode = 4'h1;
	InsTagIn = 8'h15;
#20    x_processor= 32'h0;
	y_processor= 32'h3e570a3d;
	z_processor= 32'h3ebba865;
	Opcode = 4'h2;
	InsTagIn = 8'h16;
#20    x_processor= 32'h0;
	y_processor= 32'h3e6147ae;
	z_processor= 32'h3ec49808;
	Opcode = 4'h3;
	InsTagIn = 8'h17;
#20    x_processor= 32'h0;
	y_processor= 32'h3e6b851e;
	z_processor= 32'h3ecd87ac;
	Opcode = 4'h0;
	InsTagIn = 8'h18;
#20    x_processor= 32'h0;
	y_processor= 32'h3e75c28f;
	z_processor= 32'h3ed6774f;
	Opcode = 4'h1;
	InsTagIn = 8'h19;
#20    x_processor= 32'h0;
	y_processor= 32'h3e800000;
	z_processor= 32'h3edf66f2;
	Opcode = 4'h2;
	InsTagIn = 8'h1a;
#20    x_processor= 32'h0;
	y_processor= 32'h3e851eb8;
	z_processor= 32'h3ee85696;
	Opcode = 4'h3;
	InsTagIn = 8'h1b;
#20    x_processor= 32'h0;
	y_processor= 32'h3e8a3d70;
	z_processor= 32'h3ef14639;
	Opcode = 4'h0;
	InsTagIn = 8'h1c;
#20    x_processor= 32'h0;
	y_processor= 32'h3e8f5c28;
	z_processor= 32'h3efa35dc;
	Opcode = 4'h1;
	InsTagIn = 8'h1d;
#20    x_processor= 32'h0;
	y_processor= 32'h3e947ae1;
	z_processor= 32'h3f0192c0;
	Opcode = 4'h2;
	InsTagIn = 8'h1e;
#20    x_processor= 32'h0;
	y_processor= 32'h3e999999;
	z_processor= 32'h3f060a91;
	Opcode = 4'h3;
	InsTagIn = 8'h1f;
#20    x_processor= 32'h0;
	y_processor= 32'h3e9eb851;
	z_processor= 32'h3f0a8263;
	Opcode = 4'h0;
	InsTagIn = 8'h20;
#20    x_processor= 32'h0;
	y_processor= 32'h3ea3d70a;
	z_processor= 32'h3f0efa35;
	Opcode = 4'h1;
	InsTagIn = 8'h21;
#20    x_processor= 32'h0;
	y_processor= 32'h3ea8f5c2;
	z_processor= 32'h3f137206;
	Opcode = 4'h2;
	InsTagIn = 8'h22;
#20    x_processor= 32'h3FC00000;
	y_processor= 32'h3F000000;
	z_processor= 32'h30000000;
	Opcode = 4'h5;
	InsTagIn = 8'h23;
#20    x_processor= 32'h0;
	y_processor= 32'h3eb33333;
	z_processor= 32'h3f1c61aa;
	Opcode = 4'h0;
	InsTagIn = 8'h24;
#20    x_processor= 32'h0;
	y_processor= 32'h3eb851eb;
	z_processor= 32'h3f20d97b;
	Opcode = 4'h1;
	InsTagIn = 8'h25;
#20    x_processor= 32'h0;
	y_processor= 32'h3ebd70a3;
	z_processor= 32'h3f25514d;
	Opcode = 4'h2;
	InsTagIn = 8'h26;
#20    x_processor= 32'h0;
	y_processor= 32'h3ec28f5c;
	z_processor= 32'h3f29c91f;
	Opcode = 4'h3;
	InsTagIn = 8'h27;
#20    x_processor= 32'h0;
	y_processor= 32'h3ec7ae14;
	z_processor= 32'h3f2e40f0;
	Opcode = 4'h0;
	InsTagIn = 8'h28;
#20    x_processor= 32'h0;
	y_processor= 32'h3ecccccc;
	z_processor= 32'h3f32b8c2;
	Opcode = 4'h1;
	InsTagIn = 8'h29;
//#20    x_processor= 32'h0;
//	y_processor= 32'h3ed1eb85;
//	z_processor= 32'h3f373093;
//	Opcode = 4'h2;
//	InsTagIn = 8'h2a;
#20    x_processor= 32'h00000000;
	y_processor= 32'h3FFEB852;
	z_processor= 32'h30000000;
	Opcode = 4'h9;
	InsTagIn = 8'h2a;
	
#20    x_processor= 32'h0;
	y_processor= 32'h3ed70a3d;
	z_processor= 32'h3f3ba865;
	Opcode = 4'h3;
	InsTagIn = 8'h2b;
#20    x_processor= 32'h0;
	y_processor= 32'h3edc28f5;
	z_processor= 32'h3f402037;
	Opcode = 4'h0;
	InsTagIn = 8'h2c;
#20    x_processor= 32'h0;
	y_processor= 32'h3ee147ae;
	z_processor= 32'h3f449808;
	Opcode = 4'h1;
	InsTagIn = 8'h2d;
#20    x_processor= 32'h0;
	y_processor= 32'h3ee66666;
	z_processor= 32'h3f490fda;
	Opcode = 4'h2;
	InsTagIn = 8'h2e;
#20    x_processor= 32'h0;
	y_processor= 32'h3eeb851e;
	z_processor= 32'h3f4d87ac;
	Opcode = 4'h3;
	InsTagIn = 8'h2f;
#20    x_processor= 32'h0;
	y_processor= 32'h3ef0a3d7;
	z_processor= 32'h3f51ff7d;
	Opcode = 4'h0;
	InsTagIn = 8'h30;
#20    x_processor= 32'h0;
	y_processor= 32'h3ef5c28f;
	z_processor= 32'h3f56774f;
	Opcode = 4'h1;
	InsTagIn = 8'h31;
#20    x_processor= 32'h0;
	y_processor= 32'h3efae147;
	z_processor= 32'h3f5aef21;
	Opcode = 4'h2;
	InsTagIn = 8'h32;
#20    x_processor= 32'h0;
	y_processor= 32'h3f000000;
	z_processor= 32'h3f5f66f2;
	Opcode = 4'h3;
	InsTagIn = 8'h33;
#20    x_processor= 32'h0;
	y_processor= 32'h3f028f5c;
	z_processor= 32'h3f63dec4;
	Opcode = 4'h0;
	InsTagIn = 8'h34;
#20    x_processor= 32'h0;
	y_processor= 32'h3f051eb8;
	z_processor= 32'h3f685696;
	Opcode = 4'h1;
	InsTagIn = 8'h35;
#20    x_processor= 32'h0;
	y_processor= 32'h3f07ae14;
	z_processor= 32'h3f6cce67;
	Opcode = 4'h2;
	InsTagIn = 8'h36;
#20    x_processor= 32'h0;
	y_processor= 32'h3f0a3d70;
	z_processor= 32'h3f714639;
	Opcode = 4'h3;
	InsTagIn = 8'h37;
#20    x_processor= 32'h0;
	y_processor= 32'h3f0ccccc;
	z_processor= 32'h3f75be0b;
	Opcode = 4'h0;
	InsTagIn = 8'h38;
#20    x_processor= 32'h0;
	y_processor= 32'h3f0f5c28;
	z_processor= 32'h3f7a35dc;
	Opcode = 4'h1;
	InsTagIn = 8'h39;
#20    x_processor= 32'h0;
	y_processor= 32'h3f11eb85;
	z_processor= 32'h3f7eadae;
	Opcode = 4'h2;
	InsTagIn = 8'h3a;
#20    x_processor= 32'h0;
	y_processor= 32'h3f147ae1;
	z_processor= 32'h3f8192c0;
	Opcode = 4'h3;
	InsTagIn = 8'h3b;
#20    x_processor= 32'h0;
	y_processor= 32'h3f170a3d;
	z_processor= 32'h3f83cea8;
	Opcode = 4'h0;
	InsTagIn = 8'h3c;
#20    x_processor= 32'h0;
	y_processor= 32'h3f199999;
	z_processor= 32'h3f860a91;
	Opcode = 4'h1;
	InsTagIn = 8'h3d;
#20    x_processor= 32'h0;
	y_processor= 32'h3f1c28f5;
	z_processor= 32'h3f88467a;
	Opcode = 4'h2;
	InsTagIn = 8'h3e;
#20    x_processor= 32'h0;
	y_processor= 32'h3f1eb851;
	z_processor= 32'h3f8a8263;
	Opcode = 4'h3;
	InsTagIn = 8'h3f;
#20    x_processor= 32'h0;
	y_processor= 32'h3f2147ae;
	z_processor= 32'h3f8cbe4c;
	Opcode = 4'h0;
	InsTagIn = 8'h40;
#20    x_processor= 32'h0;
	y_processor= 32'h3f23d70a;
	z_processor= 32'h3f8efa35;
	Opcode = 4'h1;
	InsTagIn = 8'h41;
#20    x_processor= 32'h0;
	y_processor= 32'h3f266666;
	z_processor= 32'h3f91361d;
	Opcode = 4'h2;
	InsTagIn = 8'h42;
#20    x_processor= 32'h0;
	y_processor= 32'h3f28f5c2;
	z_processor= 32'h3f937206;
	Opcode = 4'h3;
	InsTagIn = 8'h43;
#20    x_processor= 32'h0;
	y_processor= 32'h3f2b851e;
	z_processor= 32'h3f95adef;
	Opcode = 4'h0;
	InsTagIn = 8'h44;
#20    x_processor= 32'h0;
	y_processor= 32'h3f2e147a;
	z_processor= 32'h3f97e9d8;
	Opcode = 4'h1;
	InsTagIn = 8'h45;
#20    x_processor= 32'h0;
	y_processor= 32'h3f30a3d7;
	z_processor= 32'h3f9a25c1;
	Opcode = 4'h2;
	InsTagIn = 8'h46;
#20    x_processor= 32'h0;
	y_processor= 32'h3f333333;
	z_processor= 32'h3f9c61aa;
	Opcode = 4'h3;
	InsTagIn = 8'h47;
#20    x_processor= 32'h0;
	y_processor= 32'h3f35c28f;
	z_processor= 32'h3f9e9d92;
	Opcode = 4'h0;
	InsTagIn = 8'h48;
#20    x_processor= 32'h0;
	y_processor= 32'h3f3851eb;
	z_processor= 32'h3fa0d97b;
	Opcode = 4'h1;
	InsTagIn = 8'h49;
#20    x_processor= 32'h0;
	y_processor= 32'h3f3ae147;
	z_processor= 32'h3fa31564;
	Opcode = 4'h2;
	InsTagIn = 8'h4a;
#20    x_processor= 32'h0;
	y_processor= 32'h3f3d70a3;
	z_processor= 32'h3fa5514d;
	Opcode = 4'h3;
	InsTagIn = 8'h4b;
#20    x_processor= 32'h0;
	y_processor= 32'h3f3fffff;
	z_processor= 32'h3fa78d36;
	Opcode = 4'h0;
	InsTagIn = 8'h4c;
#20    x_processor= 32'h0;
	y_processor= 32'h3f428f5c;
	z_processor= 32'h3fa9c91f;
	Opcode = 4'h1;
	InsTagIn = 8'h4d;
#20    x_processor= 32'h0;
	y_processor= 32'h3f451eb8;
	z_processor= 32'h3fac0507;
	Opcode = 4'h2;
	InsTagIn = 8'h4e;
#20    x_processor= 32'h0;
	y_processor= 32'h3f47ae14;
	z_processor= 32'h3fae40f0;
	Opcode = 4'h3;
	InsTagIn = 8'h4f;
#20    x_processor= 32'h0;
	y_processor= 32'h3f4a3d70;
	z_processor= 32'h3fb07cd9;
	Opcode = 4'h0;
	InsTagIn = 8'h50;
#20    x_processor= 32'h0;
	y_processor= 32'h3f4ccccc;
	z_processor= 32'h3fb2b8c2;
	Opcode = 4'h1;
	InsTagIn = 8'h51;
#20    x_processor= 32'h0;
	y_processor= 32'h3f4f5c28;
	z_processor= 32'h3fb4f4ab;
	Opcode = 4'h2;
	InsTagIn = 8'h52;
#20    x_processor= 32'h0;
	y_processor= 32'h3f51eb85;
	z_processor= 32'h3fb73093;
	Opcode = 4'h3;
	InsTagIn = 8'h53;
#20    x_processor= 32'h0;
	y_processor= 32'h3f547ae1;
	z_processor= 32'h3fb96c7c;
	Opcode = 4'h0;
	InsTagIn = 8'h54;
#20    x_processor= 32'h0;
	y_processor= 32'h3f570a3d;
	z_processor= 32'h3fbba865;
	Opcode = 4'h1;
	InsTagIn = 8'h55;
#20    x_processor= 32'h0;
	y_processor= 32'h3f599999;
	z_processor= 32'h3fbde44e;
	Opcode = 4'h2;
	InsTagIn = 8'h56;
#20    x_processor= 32'h0;
	y_processor= 32'h3f5c28f5;
	z_processor= 32'h3fc02037;
	Opcode = 4'h3;
	InsTagIn = 8'h57;
#20    x_processor= 32'h0;
	y_processor= 32'h3f5eb851;
	z_processor= 32'h3fc25c20;
	Opcode = 4'h0;
	InsTagIn = 8'h58;
#20    x_processor= 32'h0;
	y_processor= 32'h3f6147ae;
	z_processor= 32'h3fc49808;
	Opcode = 4'h1;
	InsTagIn = 8'h59;
#20    x_processor= 32'h0;
	y_processor= 32'h3f63d70a;
	z_processor= 32'h3fc6d3f1;
	Opcode = 4'h2;
	InsTagIn = 8'h5a;
#20    x_processor= 32'h0;
	y_processor= 32'h3f666666;
	z_processor= 32'h3fc90fda;
	Opcode = 4'h3;
	InsTagIn = 8'h5b;
#20    x_processor= 32'h0;
	y_processor= 32'h3f68f5c2;
	z_processor= 32'h3fcb4bc3;
	Opcode = 4'h0;
	InsTagIn = 8'h5c;
#20    x_processor= 32'h0;
	y_processor= 32'h3f6b851e;
	z_processor= 32'h3fcd87ac;
	Opcode = 4'h1;
	InsTagIn = 8'h5d;
#20    x_processor= 32'h0;
	y_processor= 32'h3f6e147a;
	z_processor= 32'h3fcfc395;
	Opcode = 4'h2;
	InsTagIn = 8'h5e;
#20    x_processor= 32'h0;
	y_processor= 32'h3f70a3d7;
	z_processor= 32'h3fd1ff7d;
	Opcode = 4'h3;
	InsTagIn = 8'h5f;
#20    x_processor= 32'h0;
	y_processor= 32'h3f733333;
	z_processor= 32'h3fd43b66;
	Opcode = 4'h0;
	InsTagIn = 8'h60;
#20    x_processor= 32'h0;
	y_processor= 32'h3f75c28f;
	z_processor= 32'h3fd6774f;
	Opcode = 4'h1;
	InsTagIn = 8'h61;
#20    x_processor= 32'h0;
	y_processor= 32'h3f7851eb;
	z_processor= 32'h3fd8b338;
	Opcode = 4'h2;
	InsTagIn = 8'h62;
#20    x_processor= 32'h0;
	y_processor= 32'h3f7ae147;
	z_processor= 32'h3fdaef21;
	Opcode = 4'h3;
	InsTagIn = 8'h63;
#20    x_processor= 32'h0;
	y_processor= 32'h3f7d70a3;
	z_processor= 32'h3fdd2b0a;
	Opcode = 4'h0;
	InsTagIn = 8'h64;

end


initial begin
  f = $fopen("output1.txt");
  y = $fopen("output2.txt");
end
always@(posedge clk) begin
  repeat(20)
  begin
  $fdisplayh(f,Instruction_out);
  //$fdisplayh(y,regfile);
  end
end
always #10 clk=~clk;
always@(posedge clk)
begin
	if (OutputReady==1'b1)
	begin
	Itagregfile[i] <= Instruction_out[103:96];
	xregfile[i] <= Instruction_out[31:0];
	yregfile[i] <= Instruction_out[63:32];
	zregfile[i] <= Instruction_out[95:64];
 	i = i+1;
	end
end

always@(posedge clk)
begin
Instruction[107:100] = InsTagIn;
Instruction[99:96] = Opcode;
Instruction[31:0] = x_processor;
Instruction[63:32] = y_processor;
Instruction[95:64] = z_processor;
end
endmodule
