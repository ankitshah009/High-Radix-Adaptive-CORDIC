`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date:    14:59:40 02/21/2015 
// Design Name: 
// Module Name:    FSM_2 
// Project Name: 
// Target Devices: 
// Tool versions: 
// Description: 
//
// Dependencies: 
//
// Revision: 
// Revision 0.01 - File Created
// Additional Comments: 
//
//////////////////////////////////////////////////////////////////////////////////
module FSM_2(
    input [31:0] x_FSM1,					// x Input to FSM from Mux
    input [31:0] y_FSM1,					// y Input to FSM from Mux
    input [31:0] z_FSM1,					// z Input to FSM from Mux
    input [31:0] k_FSM1,					// k Input to FSM from Mux
	 input [31:0] theta_FSM1,
	 input [31:0] kappa_FSM1,
	 input [31:0] delta_FSM1,
    input [1:0] mode_FSM1,						// Linear: 00 Hyperbolic: 11 Circular: 01
    input operation_FSM1,							// Operation = 1 is rotation. operation = 0 is vectoring
	 input NatLogFlagout_FSM1,
	 input reset,
    input clock,
	 input [1:0] enable_LUT,				// Decides which LUT to use
	 input [7:0] address,
	 input [3:0] state_FSM2,				// State decides which part of the enabled LUT to access
	 input [7:0] InsTagFSM1Out,
	 output reg [31:0] x_FSM2,				// x_FSM1 enters FSM2
	 output reg [31:0] y_FSM2,				// y_FSM1 enters FSM2
	 output reg [31:0] z_FSM2,				// z_FSM1 enters FSM2
	 output reg [31:0] k_FSM2,				// k_FSM1 enters FSM2
    output reg [31:0] theta_FSM2,		// theta Output to ALU
    output reg [31:0] kappa_FSM2,		// kappa Output to ALU
    output reg [31:0] delta_FSM2,		// delta Output to ALU	 
	 output reg [1:0] mode_FSM2,
	 output reg operation_FSM2,
	 output reg NatLogFlagout_FSM,
	 output reg [7:0] InsTagFSMOut
    );

reg [7:0] exponent;

// Rotation LUT
reg [31:0] Rot_Theta [0:255];
reg [31:0] Rot_Delta_Cir [0:255];
reg [31:0] Rot_Delta_Hyper [0:255];
reg [31:0] Rot_Kappa_Cir [0:255];
reg [31:0] Rot_Kappa_Hyper [0:255];

// Vector LUT
reg [31:0] Vec_Theta_Cir [0:255];
reg [31:0] Vec_Theta_Hyper [0:255];
reg [31:0] Vec_Delta[0:255];
reg [31:0] Vec_Kappa_Cir [0:255];
reg [31:0] Vec_Kappa_Hyper [0:255];

// Linear Vectoring LUT
reg [31:0] LinVec_Delta [0:255];

parameter rotation  =1'b1, 
			 vectoring =1'b0;
			 
parameter mode_circular  =2'b01, 
			 mode_linear    =2'b00, 
			 mode_hyperbolic=2'b11;
			 
parameter Linear_Rotation                =  4'd0,
			 Hyperbolic_Rotation_by_1       =  4'd1,
			 Circular_Rotation_by_1         =  4'd2,
			 Rotation_with_small_theta      =  4'd3,
			 Circular_Rotation_with_table   =  4'd4,
          Hyperbolic_Rotation_with_table =  4'd5,
          Linear_Vectoring               =  4'd6,
          Hyperbolic_Vectoring_by_1      =  4'd7,
          Circular_Vectoring_by_1        =  4'd8,			 
          Vectoring_by_small_fraction    =  4'd9,
			 Circular_Vectoring_with_table  =  4'd10,
			 Hyperbolic_Vectoring_with_table=  4'd11,
			 Idle_state							  =  4'd12,
			 ConvergeRotation					  =  4'd13,
			 ConvergeVectoring				  =  4'd14;

parameter LUT_disable   = 2'b00,
			 LUT_Rotation	= 2'b01,
			 LUT_Vectoring	= 2'b10,
			 LUT_LinVec		= 2'b11;

always @ (*)
begin

	case (operation_FSM1)
	  rotation : exponent <= 8'b01111111 - z_FSM1[30:23];
	  vectoring : exponent <= y_FSM1[30:23] - x_FSM1[30:23];
	  default : exponent <= y_FSM1[30:23] - x_FSM1[30:23];
	endcase

end

always @(posedge clock)
begin


if(reset == 1'b1) begin

	// Rotation theta
	Rot_Theta[0] <=32'h3F800000;
	Rot_Theta[1] <=32'h3F800000;
	Rot_Theta[2] <=32'h3F800000;
	Rot_Theta[3] <=32'h3F800000;
	Rot_Theta[4] <=32'h3F800000;
	Rot_Theta[5] <=32'h3F800000;
	Rot_Theta[6] <=32'h3F800000;
	Rot_Theta[7] <=32'h3F800000;
	Rot_Theta[8] <=32'h3F800000;
	Rot_Theta[9] <=32'h3F800000;
	Rot_Theta[10] <=32'h3F800000;
	Rot_Theta[11] <=32'h3F800000;
	Rot_Theta[12] <=32'h3F800000;
	Rot_Theta[13] <=32'h3F800000;
	Rot_Theta[14] <=32'h3F800000;
	Rot_Theta[15] <=32'h3F800000;
	Rot_Theta[16] <=32'h3F000000;
	Rot_Theta[17] <=32'h3F080000;
	Rot_Theta[18] <=32'h3F100000;
	Rot_Theta[19] <=32'h3F180000;
	Rot_Theta[20] <=32'h3F200000;
	Rot_Theta[21] <=32'h3F280000;
	Rot_Theta[22] <=32'h3F300000;
	Rot_Theta[23] <=32'h3F380000;
	Rot_Theta[24] <=32'h3F400000;
	Rot_Theta[25] <=32'h3F480000;
	Rot_Theta[26] <=32'h3F500000;
	Rot_Theta[27] <=32'h3F580000;
	Rot_Theta[28] <=32'h3F600000;
	Rot_Theta[29] <=32'h3F680000;
	Rot_Theta[30] <=32'h3F700000;
	Rot_Theta[31] <=32'h3F780000;
	Rot_Theta[32] <=32'h3E800000;
	Rot_Theta[33] <=32'h3E880000;
	Rot_Theta[34] <=32'h3E900000;
	Rot_Theta[35] <=32'h3E980000;
	Rot_Theta[36] <=32'h3EA00000;
	Rot_Theta[37] <=32'h3EA80000;
	Rot_Theta[38] <=32'h3EB00000;
	Rot_Theta[39] <=32'h3EB80000;
	Rot_Theta[40] <=32'h3EC00000;
	Rot_Theta[41] <=32'h3EC80000;
	Rot_Theta[42] <=32'h3ED00000;
	Rot_Theta[43] <=32'h3ED80000;
	Rot_Theta[44] <=32'h3EE00000;
	Rot_Theta[45] <=32'h3EE80000;
	Rot_Theta[46] <=32'h3EF00000;
	Rot_Theta[47] <=32'h3EF80000;
	Rot_Theta[48] <=32'h3E000000;
	Rot_Theta[49] <=32'h3E080000;
	Rot_Theta[50] <=32'h3E100000;
	Rot_Theta[51] <=32'h3E180000;
	Rot_Theta[52] <=32'h3E200000;
	Rot_Theta[53] <=32'h3E280000;
	Rot_Theta[54] <=32'h3E300000;
	Rot_Theta[55] <=32'h3E380000;
	Rot_Theta[56] <=32'h3E400000;
	Rot_Theta[57] <=32'h3E480000;
	Rot_Theta[58] <=32'h3E500000;
	Rot_Theta[59] <=32'h3E580000;
	Rot_Theta[60] <=32'h3E600000;
	Rot_Theta[61] <=32'h3E680000;
	Rot_Theta[62] <=32'h3E700000;
	Rot_Theta[63] <=32'h3E780000;
	Rot_Theta[64] <=32'h3D800000;
	Rot_Theta[65] <=32'h3D880000;
	Rot_Theta[66] <=32'h3D900000;
	Rot_Theta[67] <=32'h3D980000;
	Rot_Theta[68] <=32'h3DA00000;
	Rot_Theta[69] <=32'h3DA80000;
	Rot_Theta[70] <=32'h3DB00000;
	Rot_Theta[71] <=32'h3DB80000;
	Rot_Theta[72] <=32'h3DC00000;
	Rot_Theta[73] <=32'h3DC80000;
	Rot_Theta[74] <=32'h3DD00000;
	Rot_Theta[75] <=32'h3DD80000;
	Rot_Theta[76] <=32'h3DE00000;
	Rot_Theta[77] <=32'h3DE80000;
	Rot_Theta[78] <=32'h3DF00000;
	Rot_Theta[79] <=32'h3DF80000;
	Rot_Theta[80] <=32'h3D000000;
	Rot_Theta[81] <=32'h3D080000;
	Rot_Theta[82] <=32'h3D100000;
	Rot_Theta[83] <=32'h3D180000;
	Rot_Theta[84] <=32'h3D200000;
	Rot_Theta[85] <=32'h3D280000;
	Rot_Theta[86] <=32'h3D300000;
	Rot_Theta[87] <=32'h3D380000;
	Rot_Theta[88] <=32'h3D400000;
	Rot_Theta[89] <=32'h3D480000;
	Rot_Theta[90] <=32'h3D500000;
	Rot_Theta[91] <=32'h3D580000;
	Rot_Theta[92] <=32'h3D600000;
	Rot_Theta[93] <=32'h3D680000;
	Rot_Theta[94] <=32'h3D700000;
	Rot_Theta[95] <=32'h3D780000;
	Rot_Theta[96] <=32'h3C800000;
	Rot_Theta[97] <=32'h3C880000;
	Rot_Theta[98] <=32'h3C900000;
	Rot_Theta[99] <=32'h3C980000;
	Rot_Theta[100] <=32'h3CA00000;
	Rot_Theta[101] <=32'h3CA80000;
	Rot_Theta[102] <=32'h3CB00000;
	Rot_Theta[103] <=32'h3CB80000;
	Rot_Theta[104] <=32'h3CC00000;
	Rot_Theta[105] <=32'h3CC80000;
	Rot_Theta[106] <=32'h3CD00000;
	Rot_Theta[107] <=32'h3CD80000;
	Rot_Theta[108] <=32'h3CE00000;
	Rot_Theta[109] <=32'h3CE80000;
	Rot_Theta[110] <=32'h3CF00000;
	Rot_Theta[111] <=32'h3CF80000;
	Rot_Theta[112] <=32'h3C000000;
	Rot_Theta[113] <=32'h3C080000;
	Rot_Theta[114] <=32'h3C100000;
	Rot_Theta[115] <=32'h3C180000;
	Rot_Theta[116] <=32'h3C200000;
	Rot_Theta[117] <=32'h3C280000;
	Rot_Theta[118] <=32'h3C300000;
	Rot_Theta[119] <=32'h3C380000;
	Rot_Theta[120] <=32'h3C400000;
	Rot_Theta[121] <=32'h3C480000;
	Rot_Theta[122] <=32'h3C500000;
	Rot_Theta[123] <=32'h3C580000;
	Rot_Theta[124] <=32'h3C600000;
	Rot_Theta[125] <=32'h3C680000;
	Rot_Theta[126] <=32'h3C700000;
	Rot_Theta[127] <=32'h3C780000;
	Rot_Theta[128] <=32'h3B800000;
	Rot_Theta[129] <=32'h3B880000;
	Rot_Theta[130] <=32'h3B900000;
	Rot_Theta[131] <=32'h3B980000;
	Rot_Theta[132] <=32'h3BA00000;
	Rot_Theta[133] <=32'h3BA80000;
	Rot_Theta[134] <=32'h3BB00000;
	Rot_Theta[135] <=32'h3BB80000;
	Rot_Theta[136] <=32'h3BC00000;
	Rot_Theta[137] <=32'h3BC80000;
	Rot_Theta[138] <=32'h3BD00000;
	Rot_Theta[139] <=32'h3BD80000;
	Rot_Theta[140] <=32'h3BE00000;
	Rot_Theta[141] <=32'h3BE80000;
	Rot_Theta[142] <=32'h3BF00000;
	Rot_Theta[143] <=32'h3BF80000;
	Rot_Theta[144] <=32'h3B000000;
	Rot_Theta[145] <=32'h3B080000;
	Rot_Theta[146] <=32'h3B100000;
	Rot_Theta[147] <=32'h3B180000;
	Rot_Theta[148] <=32'h3B200000;
	Rot_Theta[149] <=32'h3B280000;
	Rot_Theta[150] <=32'h3B300000;
	Rot_Theta[151] <=32'h3B380000;
	Rot_Theta[152] <=32'h3B400000;
	Rot_Theta[153] <=32'h3B480000;
	Rot_Theta[154] <=32'h3B500000;
	Rot_Theta[155] <=32'h3B580000;
	Rot_Theta[156] <=32'h3B600000;
	Rot_Theta[157] <=32'h3B680000;
	Rot_Theta[158] <=32'h3B700000;
	Rot_Theta[159] <=32'h3B780000;
	Rot_Theta[160] <=32'h3A800000;
	Rot_Theta[161] <=32'h3A880000;
	Rot_Theta[162] <=32'h3A900000;
	Rot_Theta[163] <=32'h3A980000;
	Rot_Theta[164] <=32'h3AA00000;
	Rot_Theta[165] <=32'h3AA80000;
	Rot_Theta[166] <=32'h3AB00000;
	Rot_Theta[167] <=32'h3AB80000;
	Rot_Theta[168] <=32'h3AC00000;
	Rot_Theta[169] <=32'h3AC80000;
	Rot_Theta[170] <=32'h3AD00000;
	Rot_Theta[171] <=32'h3AD80000;
	Rot_Theta[172] <=32'h3AE00000;
	Rot_Theta[173] <=32'h3AE80000;
	Rot_Theta[174] <=32'h3AF00000;
	Rot_Theta[175] <=32'h3AF80000;
	Rot_Theta[176] <=32'h3A000000;
	Rot_Theta[177] <=32'h3A080000;
	Rot_Theta[178] <=32'h3A100000;
	Rot_Theta[179] <=32'h3A180000;
	Rot_Theta[180] <=32'h3A200000;
	Rot_Theta[181] <=32'h3A280000;
	Rot_Theta[182] <=32'h3A300000;
	Rot_Theta[183] <=32'h3A380000;
	Rot_Theta[184] <=32'h3A400000;
	Rot_Theta[185] <=32'h3A480000;
	Rot_Theta[186] <=32'h3A500000;
	Rot_Theta[187] <=32'h3A580000;
	Rot_Theta[188] <=32'h3A600000;
	Rot_Theta[189] <=32'h3A680000;
	Rot_Theta[190] <=32'h3A700000;
	Rot_Theta[191] <=32'h3A780000;
	Rot_Theta[192] <=32'h39800000;
	Rot_Theta[193] <=32'h39880000;
	Rot_Theta[194] <=32'h39900000;
	Rot_Theta[195] <=32'h39980000;
	Rot_Theta[196] <=32'h39A00000;
	Rot_Theta[197] <=32'h39A80000;
	Rot_Theta[198] <=32'h39B00000;
	Rot_Theta[199] <=32'h39B80000;
	Rot_Theta[200] <=32'h39C00000;
	Rot_Theta[201] <=32'h39C80000;
	Rot_Theta[202] <=32'h39D00000;
	Rot_Theta[203] <=32'h39D80000;
	Rot_Theta[204] <=32'h39E00000;
	Rot_Theta[205] <=32'h39E80000;
	Rot_Theta[206] <=32'h39F00000;
	Rot_Theta[207] <=32'h39F80000;
	Rot_Theta[208] <=32'h39000000;
	Rot_Theta[209] <=32'h39080000;
	Rot_Theta[210] <=32'h39100000;
	Rot_Theta[211] <=32'h39180000;
	Rot_Theta[212] <=32'h39200000;
	Rot_Theta[213] <=32'h39280000;
	Rot_Theta[214] <=32'h39300000;
	Rot_Theta[215] <=32'h39380000;
	Rot_Theta[216] <=32'h39400000;
	Rot_Theta[217] <=32'h39480000;
	Rot_Theta[218] <=32'h39500000;
	Rot_Theta[219] <=32'h39580000;
	Rot_Theta[220] <=32'h39600000;
	Rot_Theta[221] <=32'h39680000;
	Rot_Theta[222] <=32'h39700000;
	Rot_Theta[223] <=32'h39780000;
	Rot_Theta[224] <=32'h38800000;
	Rot_Theta[225] <=32'h38880000;
	Rot_Theta[226] <=32'h38900000;
	Rot_Theta[227] <=32'h38980000;
	Rot_Theta[228] <=32'h38A00000;
	Rot_Theta[229] <=32'h38A80000;
	Rot_Theta[230] <=32'h38B00000;
	Rot_Theta[231] <=32'h38B80000;
	Rot_Theta[232] <=32'h38C00000;
	Rot_Theta[233] <=32'h38C80000;
	Rot_Theta[234] <=32'h38D00000;
	Rot_Theta[235] <=32'h38D80000;
	Rot_Theta[236] <=32'h38E00000;
	Rot_Theta[237] <=32'h38E80000;
	Rot_Theta[238] <=32'h38F00000;
	Rot_Theta[239] <=32'h38F80000;
	Rot_Theta[240] <=32'h38000000;
	Rot_Theta[241] <=32'h38080000;
	Rot_Theta[242] <=32'h38100000;
	Rot_Theta[243] <=32'h38180000;
	Rot_Theta[244] <=32'h38200000;
	Rot_Theta[245] <=32'h38280000;
	Rot_Theta[246] <=32'h38300000;
	Rot_Theta[247] <=32'h38380000;
	Rot_Theta[248] <=32'h38400000;
	Rot_Theta[249] <=32'h38480000;
	Rot_Theta[250] <=32'h38500000;
	Rot_Theta[251] <=32'h38580000;
	Rot_Theta[252] <=32'h38600000;
	Rot_Theta[253] <=32'h38680000;
	Rot_Theta[254] <=32'h38700000;
	Rot_Theta[255] <=32'h38780000;

	// Rotation delta for circular mode
	Rot_Delta_Cir[0] <=32'h3FC75922;
	Rot_Delta_Cir[1] <=32'h3FC75922;
	Rot_Delta_Cir[2] <=32'h3FC75922;
	Rot_Delta_Cir[3] <=32'h3FC75922;
	Rot_Delta_Cir[4] <=32'h3FC75922;
	Rot_Delta_Cir[5] <=32'h3FC75922;
	Rot_Delta_Cir[6] <=32'h3FC75922;
	Rot_Delta_Cir[7] <=32'h3FC75922;
	Rot_Delta_Cir[8] <=32'h3FC75922;
	Rot_Delta_Cir[9] <=32'h3FC75922;
	Rot_Delta_Cir[10] <=32'h3FC75922;
	Rot_Delta_Cir[11] <=32'h3FC75922;
	Rot_Delta_Cir[12] <=32'h3FC75922;
	Rot_Delta_Cir[13] <=32'h3FC75922;
	Rot_Delta_Cir[14] <=32'h3FC75922;
	Rot_Delta_Cir[15] <=32'h3FC75922;
	Rot_Delta_Cir[16] <=32'h3F0BDA7A;
	Rot_Delta_Cir[17] <=32'h3F166CC7;
	Rot_Delta_Cir[18] <=32'h3F21645D;
	Rot_Delta_Cir[19] <=32'h3F2CCCD4;
	Rot_Delta_Cir[20] <=32'h3F38B334;
	Rot_Delta_Cir[21] <=32'h3F452629;
	Rot_Delta_Cir[22] <=32'h3F523659;
	Rot_Delta_Cir[23] <=32'h3F5FF6BE;
	Rot_Delta_Cir[24] <=32'h3F6E7D1B;
	Rot_Delta_Cir[25] <=32'h3F7DE288;
	Rot_Delta_Cir[26] <=32'h3F872215;
	Rot_Delta_Cir[27] <=32'h3F8FE205;
	Rot_Delta_Cir[28] <=32'h3F99451C;
	Rot_Delta_Cir[29] <=32'h3FA36319;
	Rot_Delta_Cir[30] <=32'h3FAE585F;
	Rot_Delta_Cir[31] <=32'h3FBA4729;
	Rot_Delta_Cir[32] <=32'h3E82BC2D;
	Rot_Delta_Cir[33] <=32'h3E8B4A9F;
	Rot_Delta_Cir[34] <=32'h3E93EBC5;
	Rot_Delta_Cir[35] <=32'h3E9CA0F5;
	Rot_Delta_Cir[36] <=32'h3EA56B8F;
	Rot_Delta_Cir[37] <=32'h3EAE4D00;
	Rot_Delta_Cir[38] <=32'h3EB746C2;
	Rot_Delta_Cir[39] <=32'h3EC05A5E;
	Rot_Delta_Cir[40] <=32'h3EC9896C;
	Rot_Delta_Cir[41] <=32'h3ED2D593;
	Rot_Delta_Cir[42] <=32'h3EDC408F;
	Rot_Delta_Cir[43] <=32'h3EE5CC2C;
	Rot_Delta_Cir[44] <=32'h3EEF7A4F;
	Rot_Delta_Cir[45] <=32'h3EF94CEF;
	Rot_Delta_Cir[46] <=32'h3F01A30F;
	Rot_Delta_Cir[47] <=32'h3F06B404;
	Rot_Delta_Cir[48] <=32'h3E00ABBD;
	Rot_Delta_Cir[49] <=32'h3E08CE29;
	Rot_Delta_Cir[50] <=32'h3E10F4F0;
	Rot_Delta_Cir[51] <=32'h3E192055;
	Rot_Delta_Cir[52] <=32'h3E21509E;
	Rot_Delta_Cir[53] <=32'h3E298613;
	Rot_Delta_Cir[54] <=32'h3E31C0F9;
	Rot_Delta_Cir[55] <=32'h3E3A0197;
	Rot_Delta_Cir[56] <=32'h3E424837;
	Rot_Delta_Cir[57] <=32'h3E4A9521;
	Rot_Delta_Cir[58] <=32'h3E52E89F;
	Rot_Delta_Cir[59] <=32'h3E5B42FD;
	Rot_Delta_Cir[60] <=32'h3E63A485;
	Rot_Delta_Cir[61] <=32'h3E6C0D84;
	Rot_Delta_Cir[62] <=32'h3E747E48;
	Rot_Delta_Cir[63] <=32'h3E7CF71F;
	Rot_Delta_Cir[64] <=32'h3D802ABB;
	Rot_Delta_Cir[65] <=32'h3D883344;
	Rot_Delta_Cir[66] <=32'h3D903CDE;
	Rot_Delta_Cir[67] <=32'h3D98479B;
	Rot_Delta_Cir[68] <=32'h3DA05389;
	Rot_Delta_Cir[69] <=32'h3DA860BA;
	Rot_Delta_Cir[70] <=32'h3DB06F3E;
	Rot_Delta_Cir[71] <=32'h3DB87F26;
	Rot_Delta_Cir[72] <=32'h3DC09082;
	Rot_Delta_Cir[73] <=32'h3DC8A362;
	Rot_Delta_Cir[74] <=32'h3DD0B7D7;
	Rot_Delta_Cir[75] <=32'h3DD8CDF2;
	Rot_Delta_Cir[76] <=32'h3DE0E5C4;
	Rot_Delta_Cir[77] <=32'h3DE8FF5C;
	Rot_Delta_Cir[78] <=32'h3DF11ACD;
	Rot_Delta_Cir[79] <=32'h3DF93827;
	Rot_Delta_Cir[80] <=32'h3D000AAB;
	Rot_Delta_Cir[81] <=32'h3D080CCC;
	Rot_Delta_Cir[82] <=32'h3D100F31;
	Rot_Delta_Cir[83] <=32'h3D1811DF;
	Rot_Delta_Cir[84] <=32'h3D2014D8;
	Rot_Delta_Cir[85] <=32'h3D281822;
	Rot_Delta_Cir[86] <=32'h3D301BBF;
	Rot_Delta_Cir[87] <=32'h3D381FB5;
	Rot_Delta_Cir[88] <=32'h3D402408;
	Rot_Delta_Cir[89] <=32'h3D4828BA;
	Rot_Delta_Cir[90] <=32'h3D502DD1;
	Rot_Delta_Cir[91] <=32'h3D583350;
	Rot_Delta_Cir[92] <=32'h3D60393C;
	Rot_Delta_Cir[93] <=32'h3D683F98;
	Rot_Delta_Cir[94] <=32'h3D704668;
	Rot_Delta_Cir[95] <=32'h3D784DB1;
	Rot_Delta_Cir[96] <=32'h3C8002AA;
	Rot_Delta_Cir[97] <=32'h3C880332;
	Rot_Delta_Cir[98] <=32'h3C9003CC;
	Rot_Delta_Cir[99] <=32'h3C980477;
	Rot_Delta_Cir[100] <=32'h3CA00535;
	Rot_Delta_Cir[101] <=32'h3CA80607;
	Rot_Delta_Cir[102] <=32'h3CB006EE;
	Rot_Delta_Cir[103] <=32'h3CB807EC;
	Rot_Delta_Cir[104] <=32'h3CC00900;
	Rot_Delta_Cir[105] <=32'h3CC80A2C;
	Rot_Delta_Cir[106] <=32'h3CD00B72;
	Rot_Delta_Cir[107] <=32'h3CD80CD1;
	Rot_Delta_Cir[108] <=32'h3CE00E4B;
	Rot_Delta_Cir[109] <=32'h3CE80FE2;
	Rot_Delta_Cir[110] <=32'h3CF01195;
	Rot_Delta_Cir[111] <=32'h3CF81366;
	Rot_Delta_Cir[112] <=32'h3C0000AA;
	Rot_Delta_Cir[113] <=32'h3C0800CC;
	Rot_Delta_Cir[114] <=32'h3C1000F3;
	Rot_Delta_Cir[115] <=32'h3C18011D;
	Rot_Delta_Cir[116] <=32'h3C20014D;
	Rot_Delta_Cir[117] <=32'h3C280181;
	Rot_Delta_Cir[118] <=32'h3C3001BB;
	Rot_Delta_Cir[119] <=32'h3C3801FA;
	Rot_Delta_Cir[120] <=32'h3C400240;
	Rot_Delta_Cir[121] <=32'h3C48028B;
	Rot_Delta_Cir[122] <=32'h3C5002DC;
	Rot_Delta_Cir[123] <=32'h3C580334;
	Rot_Delta_Cir[124] <=32'h3C600392;
	Rot_Delta_Cir[125] <=32'h3C6803F8;
	Rot_Delta_Cir[126] <=32'h3C700465;
	Rot_Delta_Cir[127] <=32'h3C7804D9;
	Rot_Delta_Cir[128] <=32'h3B80002A;
	Rot_Delta_Cir[129] <=32'h3B880033;
	Rot_Delta_Cir[130] <=32'h3B90003C;
	Rot_Delta_Cir[131] <=32'h3B980047;
	Rot_Delta_Cir[132] <=32'h3BA00053;
	Rot_Delta_Cir[133] <=32'h3BA80060;
	Rot_Delta_Cir[134] <=32'h3BB0006E;
	Rot_Delta_Cir[135] <=32'h3BB8007E;
	Rot_Delta_Cir[136] <=32'h3BC00090;
	Rot_Delta_Cir[137] <=32'h3BC800A2;
	Rot_Delta_Cir[138] <=32'h3BD000B7;
	Rot_Delta_Cir[139] <=32'h3BD800CD;
	Rot_Delta_Cir[140] <=32'h3BE000E4;
	Rot_Delta_Cir[141] <=32'h3BE800FE;
	Rot_Delta_Cir[142] <=32'h3BF00119;
	Rot_Delta_Cir[143] <=32'h3BF80136;
	Rot_Delta_Cir[144] <=32'h3B00000A;
	Rot_Delta_Cir[145] <=32'h3B08000C;
	Rot_Delta_Cir[146] <=32'h3B10000F;
	Rot_Delta_Cir[147] <=32'h3B180011;
	Rot_Delta_Cir[148] <=32'h3B200014;
	Rot_Delta_Cir[149] <=32'h3B280018;
	Rot_Delta_Cir[150] <=32'h3B30001B;
	Rot_Delta_Cir[151] <=32'h3B38001F;
	Rot_Delta_Cir[152] <=32'h3B400024;
	Rot_Delta_Cir[153] <=32'h3B480028;
	Rot_Delta_Cir[154] <=32'h3B50002D;
	Rot_Delta_Cir[155] <=32'h3B580033;
	Rot_Delta_Cir[156] <=32'h3B600039;
	Rot_Delta_Cir[157] <=32'h3B68003F;
	Rot_Delta_Cir[158] <=32'h3B700046;
	Rot_Delta_Cir[159] <=32'h3B78004D;
	Rot_Delta_Cir[160] <=32'h3A800002;
	Rot_Delta_Cir[161] <=32'h3A880003;
	Rot_Delta_Cir[162] <=32'h3A900003;
	Rot_Delta_Cir[163] <=32'h3A980004;
	Rot_Delta_Cir[164] <=32'h3AA00005;
	Rot_Delta_Cir[165] <=32'h3AA80006;
	Rot_Delta_Cir[166] <=32'h3AB00006;
	Rot_Delta_Cir[167] <=32'h3AB80007;
	Rot_Delta_Cir[168] <=32'h3AC00009;
	Rot_Delta_Cir[169] <=32'h3AC8000A;
	Rot_Delta_Cir[170] <=32'h3AD0000B;
	Rot_Delta_Cir[171] <=32'h3AD8000C;
	Rot_Delta_Cir[172] <=32'h3AE0000E;
	Rot_Delta_Cir[173] <=32'h3AE8000F;
	Rot_Delta_Cir[174] <=32'h3AF00011;
	Rot_Delta_Cir[175] <=32'h3AF80013;
	Rot_Delta_Cir[176] <=32'h3A000000;
	Rot_Delta_Cir[177] <=32'h3A080000;
	Rot_Delta_Cir[178] <=32'h3A100000;
	Rot_Delta_Cir[179] <=32'h3A180001;
	Rot_Delta_Cir[180] <=32'h3A200001;
	Rot_Delta_Cir[181] <=32'h3A280001;
	Rot_Delta_Cir[182] <=32'h3A300001;
	Rot_Delta_Cir[183] <=32'h3A380001;
	Rot_Delta_Cir[184] <=32'h3A400002;
	Rot_Delta_Cir[185] <=32'h3A480002;
	Rot_Delta_Cir[186] <=32'h3A500002;
	Rot_Delta_Cir[187] <=32'h3A580003;
	Rot_Delta_Cir[188] <=32'h3A600003;
	Rot_Delta_Cir[189] <=32'h3A680003;
	Rot_Delta_Cir[190] <=32'h3A700004;
	Rot_Delta_Cir[191] <=32'h3A780004;
	Rot_Delta_Cir[192] <=32'h39800000;
	Rot_Delta_Cir[193] <=32'h39880000;
	Rot_Delta_Cir[194] <=32'h39900000;
	Rot_Delta_Cir[195] <=32'h39980000;
	Rot_Delta_Cir[196] <=32'h39A00000;
	Rot_Delta_Cir[197] <=32'h39A80000;
	Rot_Delta_Cir[198] <=32'h39B00000;
	Rot_Delta_Cir[199] <=32'h39B80000;
	Rot_Delta_Cir[200] <=32'h39C00000;
	Rot_Delta_Cir[201] <=32'h39C80000;
	Rot_Delta_Cir[202] <=32'h39D00000;
	Rot_Delta_Cir[203] <=32'h39D80000;
	Rot_Delta_Cir[204] <=32'h39E00000;
	Rot_Delta_Cir[205] <=32'h39E80000;
	Rot_Delta_Cir[206] <=32'h39F00001;
	Rot_Delta_Cir[207] <=32'h39F80001;
	Rot_Delta_Cir[208] <=32'h39000000;
	Rot_Delta_Cir[209] <=32'h39080000;
	Rot_Delta_Cir[210] <=32'h39100000;
	Rot_Delta_Cir[211] <=32'h39180000;
	Rot_Delta_Cir[212] <=32'h39200000;
	Rot_Delta_Cir[213] <=32'h39280000;
	Rot_Delta_Cir[214] <=32'h39300000;
	Rot_Delta_Cir[215] <=32'h39380000;
	Rot_Delta_Cir[216] <=32'h39400000;
	Rot_Delta_Cir[217] <=32'h39480000;
	Rot_Delta_Cir[218] <=32'h39500000;
	Rot_Delta_Cir[219] <=32'h39580000;
	Rot_Delta_Cir[220] <=32'h39600000;
	Rot_Delta_Cir[221] <=32'h39680000;
	Rot_Delta_Cir[222] <=32'h39700000;
	Rot_Delta_Cir[223] <=32'h39780000;
	Rot_Delta_Cir[224] <=32'h38800000;
	Rot_Delta_Cir[225] <=32'h38880000;
	Rot_Delta_Cir[226] <=32'h38900000;
	Rot_Delta_Cir[227] <=32'h38980000;
	Rot_Delta_Cir[228] <=32'h38A00000;
	Rot_Delta_Cir[229] <=32'h38A80000;
	Rot_Delta_Cir[230] <=32'h38B00000;
	Rot_Delta_Cir[231] <=32'h38B80000;
	Rot_Delta_Cir[232] <=32'h38C00000;
	Rot_Delta_Cir[233] <=32'h38C80000;
	Rot_Delta_Cir[234] <=32'h38D00000;
	Rot_Delta_Cir[235] <=32'h38D80000;
	Rot_Delta_Cir[236] <=32'h38E00000;
	Rot_Delta_Cir[237] <=32'h38E80000;
	Rot_Delta_Cir[238] <=32'h38F00000;
	Rot_Delta_Cir[239] <=32'h38F80000;
	Rot_Delta_Cir[240] <=32'h38000000;
	Rot_Delta_Cir[241] <=32'h38080000;
	Rot_Delta_Cir[242] <=32'h38100000;
	Rot_Delta_Cir[243] <=32'h38180000;
	Rot_Delta_Cir[244] <=32'h38200000;
	Rot_Delta_Cir[245] <=32'h38280000;
	Rot_Delta_Cir[246] <=32'h38300000;
	Rot_Delta_Cir[247] <=32'h38380000;
	Rot_Delta_Cir[248] <=32'h38400000;
	Rot_Delta_Cir[249] <=32'h38480000;
	Rot_Delta_Cir[250] <=32'h38500000;
	Rot_Delta_Cir[251] <=32'h38580000;
	Rot_Delta_Cir[252] <=32'h38600000;
	Rot_Delta_Cir[253] <=32'h38680000;
	Rot_Delta_Cir[254] <=32'h38700000;
	Rot_Delta_Cir[255] <=32'h38780000;

	// Rotation Delta Hyperbolic mode
	Rot_Delta_Hyper[0] <=32'h3F42F7D5;
	Rot_Delta_Hyper[1] <=32'h3F495FD9;
	Rot_Delta_Hyper[2] <=32'h3F4F2E5A;
	Rot_Delta_Hyper[3] <=32'h3F546DE5;
	Rot_Delta_Hyper[4] <=32'h3F59291D;
	Rot_Delta_Hyper[5] <=32'h3F5D6A85;
	Rot_Delta_Hyper[6] <=32'h3F613C52;
	Rot_Delta_Hyper[7] <=32'h3F64A851;
	Rot_Delta_Hyper[8] <=32'h3F67B7CB;
	Rot_Delta_Hyper[9] <=32'h3F6A737A;
	Rot_Delta_Hyper[10] <=32'h3F6CE37D;
	Rot_Delta_Hyper[11] <=32'h3F6F0F5A;
	Rot_Delta_Hyper[12] <=32'h3F70FDFC;
	Rot_Delta_Hyper[13] <=32'h3F72B5B7;
	Rot_Delta_Hyper[14] <=32'h3F743C4F;
	Rot_Delta_Hyper[15] <=32'h3F7596FF;
	Rot_Delta_Hyper[16] <=32'h3EEC9A9E;
	Rot_Delta_Hyper[17] <=32'h3EF90108;
	Rot_Delta_Hyper[18] <=32'h3F028437;
	Rot_Delta_Hyper[19] <=32'h3F0857A3;
	Rot_Delta_Hyper[20] <=32'h3F0DFA3F;
	Rot_Delta_Hyper[21] <=32'h3F136BB7;
	Rot_Delta_Hyper[22] <=32'h3F18ABEF;
	Rot_Delta_Hyper[23] <=32'h3F1DBAFC;
	Rot_Delta_Hyper[24] <=32'h3F22991F;
	Rot_Delta_Hyper[25] <=32'h3F2746C4;
	Rot_Delta_Hyper[26] <=32'h3F2BC47F;
	Rot_Delta_Hyper[27] <=32'h3F301304;
	Rot_Delta_Hyper[28] <=32'h3F343328;
	Rot_Delta_Hyper[29] <=32'h3F3825D8;
	Rot_Delta_Hyper[30] <=32'h3F3BEC1C;
	Rot_Delta_Hyper[31] <=32'h3F3F870D;
	Rot_Delta_Hyper[32] <=32'h3E7ACBF5;
	Rot_Delta_Hyper[33] <=32'h3E84E3A2;
	Rot_Delta_Hyper[34] <=32'h3E8C51CC;
	Rot_Delta_Hyper[35] <=32'h3E93AFBF;
	Rot_Delta_Hyper[36] <=32'h3E9AFCC5;
	Rot_Delta_Hyper[37] <=32'h3EA23832;
	Rot_Delta_Hyper[38] <=32'h3EA96162;
	Rot_Delta_Hyper[39] <=32'h3EB077B8;
	Rot_Delta_Hyper[40] <=32'h3EB77A9E;
	Rot_Delta_Hyper[41] <=32'h3EBE6988;
	Rot_Delta_Hyper[42] <=32'h3EC543F0;
	Rot_Delta_Hyper[43] <=32'h3ECC0959;
	Rot_Delta_Hyper[44] <=32'h3ED2B94F;
	Rot_Delta_Hyper[45] <=32'h3ED95364;
	Rot_Delta_Hyper[46] <=32'h3EDFD735;
	Rot_Delta_Hyper[47] <=32'h3EE64464;
	Rot_Delta_Hyper[48] <=32'h3DFEACC9;
	Rot_Delta_Hyper[49] <=32'h3E0734B9;
	Rot_Delta_Hyper[50] <=32'h3E0F0EE8;
	Rot_Delta_Hyper[51] <=32'h3E16E4B4;
	Rot_Delta_Hyper[52] <=32'h3E1EB5E3;
	Rot_Delta_Hyper[53] <=32'h3E26823C;
	Rot_Delta_Hyper[54] <=32'h3E2E4983;
	Rot_Delta_Hyper[55] <=32'h3E360B81;
	Rot_Delta_Hyper[56] <=32'h3E3DC7FC;
	Rot_Delta_Hyper[57] <=32'h3E457EBD;
	Rot_Delta_Hyper[58] <=32'h3E4D2F8D;
	Rot_Delta_Hyper[59] <=32'h3E54DA36;
	Rot_Delta_Hyper[60] <=32'h3E5C7E82;
	Rot_Delta_Hyper[61] <=32'h3E641C3B;
	Rot_Delta_Hyper[62] <=32'h3E6BB32E;
	Rot_Delta_Hyper[63] <=32'h3E734327;
	Rot_Delta_Hyper[64] <=32'h3D7FAACC;
	Rot_Delta_Hyper[65] <=32'h3D87CCE9;
	Rot_Delta_Hyper[66] <=32'h3D8FC35E;
	Rot_Delta_Hyper[67] <=32'h3D97B8B5;
	Rot_Delta_Hyper[68] <=32'h3D9FACDE;
	Rot_Delta_Hyper[69] <=32'h3DA79FCA;
	Rot_Delta_Hyper[70] <=32'h3DAF9168;
	Rot_Delta_Hyper[71] <=32'h3DB781AB;
	Rot_Delta_Hyper[72] <=32'h3DBF7081;
	Rot_Delta_Hyper[73] <=32'h3DC75DDB;
	Rot_Delta_Hyper[74] <=32'h3DCF49AB;
	Rot_Delta_Hyper[75] <=32'h3DD733E0;
	Rot_Delta_Hyper[76] <=32'h3DDF1C6C;
	Rot_Delta_Hyper[77] <=32'h3DE7033E;
	Rot_Delta_Hyper[78] <=32'h3DEEE849;
	Rot_Delta_Hyper[79] <=32'h3DF6CB7C;
	Rot_Delta_Hyper[80] <=32'h3CFFEAAC;
	Rot_Delta_Hyper[81] <=32'h3D07F336;
	Rot_Delta_Hyper[82] <=32'h3D0FF0D1;
	Rot_Delta_Hyper[83] <=32'h3D17EE25;
	Rot_Delta_Hyper[84] <=32'h3D1FEB2D;
	Rot_Delta_Hyper[85] <=32'h3D27E7E6;
	Rot_Delta_Hyper[86] <=32'h3D2FE44A;
	Rot_Delta_Hyper[87] <=32'h3D37E057;
	Rot_Delta_Hyper[88] <=32'h3D3FDC08;
	Rot_Delta_Hyper[89] <=32'h3D47D759;
	Rot_Delta_Hyper[90] <=32'h3D4FD246;
	Rot_Delta_Hyper[91] <=32'h3D57CCCC;
	Rot_Delta_Hyper[92] <=32'h3D5FC6E6;
	Rot_Delta_Hyper[93] <=32'h3D67C091;
	Rot_Delta_Hyper[94] <=32'h3D6FB9C8;
	Rot_Delta_Hyper[95] <=32'h3D77B288;
	Rot_Delta_Hyper[96] <=32'h3C7FFAAA;
	Rot_Delta_Hyper[97] <=32'h3C87FCCD;
	Rot_Delta_Hyper[98] <=32'h3C8FFC34;
	Rot_Delta_Hyper[99] <=32'h3C97FB88;
	Rot_Delta_Hyper[100] <=32'h3C9FFACA;
	Rot_Delta_Hyper[101] <=32'h3CA7F9F8;
	Rot_Delta_Hyper[102] <=32'h3CAFF911;
	Rot_Delta_Hyper[103] <=32'h3CB7F814;
	Rot_Delta_Hyper[104] <=32'h3CBFF700;
	Rot_Delta_Hyper[105] <=32'h3CC7F5D4;
	Rot_Delta_Hyper[106] <=32'h3CCFF48F;
	Rot_Delta_Hyper[107] <=32'h3CD7F330;
	Rot_Delta_Hyper[108] <=32'h3CDFF1B6;
	Rot_Delta_Hyper[109] <=32'h3CE7F020;
	Rot_Delta_Hyper[110] <=32'h3CEFEE6D;
	Rot_Delta_Hyper[111] <=32'h3CF7EC9C;
	Rot_Delta_Hyper[112] <=32'h3BFFFEAA;
	Rot_Delta_Hyper[113] <=32'h3C07FF33;
	Rot_Delta_Hyper[114] <=32'h3C0FFF0D;
	Rot_Delta_Hyper[115] <=32'h3C17FEE2;
	Rot_Delta_Hyper[116] <=32'h3C1FFEB2;
	Rot_Delta_Hyper[117] <=32'h3C27FE7E;
	Rot_Delta_Hyper[118] <=32'h3C2FFE44;
	Rot_Delta_Hyper[119] <=32'h3C37FE05;
	Rot_Delta_Hyper[120] <=32'h3C3FFDC0;
	Rot_Delta_Hyper[121] <=32'h3C47FD74;
	Rot_Delta_Hyper[122] <=32'h3C4FFD23;
	Rot_Delta_Hyper[123] <=32'h3C57FCCB;
	Rot_Delta_Hyper[124] <=32'h3C5FFC6D;
	Rot_Delta_Hyper[125] <=32'h3C67FC07;
	Rot_Delta_Hyper[126] <=32'h3C6FFB9B;
	Rot_Delta_Hyper[127] <=32'h3C77FB26;
	Rot_Delta_Hyper[128] <=32'h3B7FFFAA;
	Rot_Delta_Hyper[129] <=32'h3B87FFCC;
	Rot_Delta_Hyper[130] <=32'h3B8FFFC3;
	Rot_Delta_Hyper[131] <=32'h3B97FFB8;
	Rot_Delta_Hyper[132] <=32'h3B9FFFAC;
	Rot_Delta_Hyper[133] <=32'h3BA7FF9F;
	Rot_Delta_Hyper[134] <=32'h3BAFFF91;
	Rot_Delta_Hyper[135] <=32'h3BB7FF81;
	Rot_Delta_Hyper[136] <=32'h3BBFFF70;
	Rot_Delta_Hyper[137] <=32'h3BC7FF5D;
	Rot_Delta_Hyper[138] <=32'h3BCFFF48;
	Rot_Delta_Hyper[139] <=32'h3BD7FF32;
	Rot_Delta_Hyper[140] <=32'h3BDFFF1B;
	Rot_Delta_Hyper[141] <=32'h3BE7FF01;
	Rot_Delta_Hyper[142] <=32'h3BEFFEE6;
	Rot_Delta_Hyper[143] <=32'h3BF7FEC9;
	Rot_Delta_Hyper[144] <=32'h3AFFFFEA;
	Rot_Delta_Hyper[145] <=32'h3B07FFF3;
	Rot_Delta_Hyper[146] <=32'h3B0FFFF0;
	Rot_Delta_Hyper[147] <=32'h3B17FFEE;
	Rot_Delta_Hyper[148] <=32'h3B1FFFEB;
	Rot_Delta_Hyper[149] <=32'h3B27FFE7;
	Rot_Delta_Hyper[150] <=32'h3B2FFFE4;
	Rot_Delta_Hyper[151] <=32'h3B37FFE0;
	Rot_Delta_Hyper[152] <=32'h3B3FFFDC;
	Rot_Delta_Hyper[153] <=32'h3B47FFD7;
	Rot_Delta_Hyper[154] <=32'h3B4FFFD2;
	Rot_Delta_Hyper[155] <=32'h3B57FFCC;
	Rot_Delta_Hyper[156] <=32'h3B5FFFC6;
	Rot_Delta_Hyper[157] <=32'h3B67FFC0;
	Rot_Delta_Hyper[158] <=32'h3B6FFFB9;
	Rot_Delta_Hyper[159] <=32'h3B77FFB2;
	Rot_Delta_Hyper[160] <=32'h3A7FFFFA;
	Rot_Delta_Hyper[161] <=32'h3A87FFFC;
	Rot_Delta_Hyper[162] <=32'h3A8FFFFC;
	Rot_Delta_Hyper[163] <=32'h3A97FFFB;
	Rot_Delta_Hyper[164] <=32'h3A9FFFFA;
	Rot_Delta_Hyper[165] <=32'h3AA7FFF9;
	Rot_Delta_Hyper[166] <=32'h3AAFFFF9;
	Rot_Delta_Hyper[167] <=32'h3AB7FFF8;
	Rot_Delta_Hyper[168] <=32'h3ABFFFF7;
	Rot_Delta_Hyper[169] <=32'h3AC7FFF5;
	Rot_Delta_Hyper[170] <=32'h3ACFFFF4;
	Rot_Delta_Hyper[171] <=32'h3AD7FFF3;
	Rot_Delta_Hyper[172] <=32'h3ADFFFF1;
	Rot_Delta_Hyper[173] <=32'h3AE7FFF0;
	Rot_Delta_Hyper[174] <=32'h3AEFFFEE;
	Rot_Delta_Hyper[175] <=32'h3AF7FFEC;
	Rot_Delta_Hyper[176] <=32'h39FFFFFE;
	Rot_Delta_Hyper[177] <=32'h3A07FFFF;
	Rot_Delta_Hyper[178] <=32'h3A0FFFFF;
	Rot_Delta_Hyper[179] <=32'h3A17FFFE;
	Rot_Delta_Hyper[180] <=32'h3A1FFFFE;
	Rot_Delta_Hyper[181] <=32'h3A27FFFE;
	Rot_Delta_Hyper[182] <=32'h3A2FFFFE;
	Rot_Delta_Hyper[183] <=32'h3A37FFFE;
	Rot_Delta_Hyper[184] <=32'h3A3FFFFD;
	Rot_Delta_Hyper[185] <=32'h3A47FFFD;
	Rot_Delta_Hyper[186] <=32'h3A4FFFFD;
	Rot_Delta_Hyper[187] <=32'h3A57FFFC;
	Rot_Delta_Hyper[188] <=32'h3A5FFFFC;
	Rot_Delta_Hyper[189] <=32'h3A67FFFC;
	Rot_Delta_Hyper[190] <=32'h3A6FFFFB;
	Rot_Delta_Hyper[191] <=32'h3A77FFFB;
	Rot_Delta_Hyper[192] <=32'h397FFFFF;
	Rot_Delta_Hyper[193] <=32'h3987FFFF;
	Rot_Delta_Hyper[194] <=32'h398FFFFF;
	Rot_Delta_Hyper[195] <=32'h3997FFFF;
	Rot_Delta_Hyper[196] <=32'h399FFFFF;
	Rot_Delta_Hyper[197] <=32'h39A7FFFF;
	Rot_Delta_Hyper[198] <=32'h39AFFFFF;
	Rot_Delta_Hyper[199] <=32'h39B7FFFF;
	Rot_Delta_Hyper[200] <=32'h39BFFFFF;
	Rot_Delta_Hyper[201] <=32'h39C7FFFF;
	Rot_Delta_Hyper[202] <=32'h39CFFFFF;
	Rot_Delta_Hyper[203] <=32'h39D7FFFF;
	Rot_Delta_Hyper[204] <=32'h39DFFFFF;
	Rot_Delta_Hyper[205] <=32'h39E7FFFF;
	Rot_Delta_Hyper[206] <=32'h39EFFFFE;
	Rot_Delta_Hyper[207] <=32'h39F7FFFE;
	Rot_Delta_Hyper[208] <=32'h38FFFFFF;
	Rot_Delta_Hyper[209] <=32'h3907FFFF;
	Rot_Delta_Hyper[210] <=32'h390FFFFF;
	Rot_Delta_Hyper[211] <=32'h3917FFFF;
	Rot_Delta_Hyper[212] <=32'h391FFFFF;
	Rot_Delta_Hyper[213] <=32'h3927FFFF;
	Rot_Delta_Hyper[214] <=32'h392FFFFF;
	Rot_Delta_Hyper[215] <=32'h3937FFFF;
	Rot_Delta_Hyper[216] <=32'h393FFFFF;
	Rot_Delta_Hyper[217] <=32'h3947FFFF;
	Rot_Delta_Hyper[218] <=32'h394FFFFF;
	Rot_Delta_Hyper[219] <=32'h3957FFFF;
	Rot_Delta_Hyper[220] <=32'h395FFFFF;
	Rot_Delta_Hyper[221] <=32'h3967FFFF;
	Rot_Delta_Hyper[222] <=32'h396FFFFF;
	Rot_Delta_Hyper[223] <=32'h3977FFFF;
	Rot_Delta_Hyper[224] <=32'h387FFFFF;
	Rot_Delta_Hyper[225] <=32'h3887FFFF;
	Rot_Delta_Hyper[226] <=32'h388FFFFF;
	Rot_Delta_Hyper[227] <=32'h3897FFFF;
	Rot_Delta_Hyper[228] <=32'h389FFFFF;
	Rot_Delta_Hyper[229] <=32'h38A7FFFF;
	Rot_Delta_Hyper[230] <=32'h38AFFFFF;
	Rot_Delta_Hyper[231] <=32'h38B7FFFF;
	Rot_Delta_Hyper[232] <=32'h38BFFFFF;
	Rot_Delta_Hyper[233] <=32'h38C7FFFF;
	Rot_Delta_Hyper[234] <=32'h38CFFFFF;
	Rot_Delta_Hyper[235] <=32'h38D7FFFF;
	Rot_Delta_Hyper[236] <=32'h38DFFFFF;
	Rot_Delta_Hyper[237] <=32'h38E7FFFF;
	Rot_Delta_Hyper[238] <=32'h38EFFFFF;
	Rot_Delta_Hyper[239] <=32'h38F7FFFF;
	Rot_Delta_Hyper[240] <=32'h37FFFFFF;
	Rot_Delta_Hyper[241] <=32'h3807FFFF;
	Rot_Delta_Hyper[242] <=32'h380FFFFF;
	Rot_Delta_Hyper[243] <=32'h3817FFFF;
	Rot_Delta_Hyper[244] <=32'h381FFFFF;
	Rot_Delta_Hyper[245] <=32'h3827FFFF;
	Rot_Delta_Hyper[246] <=32'h382FFFFF;
	Rot_Delta_Hyper[247] <=32'h3837FFFF;
	Rot_Delta_Hyper[248] <=32'h383FFFFF;
	Rot_Delta_Hyper[249] <=32'h3847FFFF;
	Rot_Delta_Hyper[250] <=32'h384FFFFF;
	Rot_Delta_Hyper[251] <=32'h3857FFFF;
	Rot_Delta_Hyper[252] <=32'h385FFFFF;
	Rot_Delta_Hyper[253] <=32'h3867FFFF;
	Rot_Delta_Hyper[254] <=32'h386FFFFF;
	Rot_Delta_Hyper[255] <=32'h3877FFFF;
	
	// Rotation Kappa Circular
	Rot_Kappa_Cir[0] <=32'h3F0A5142;
	Rot_Kappa_Cir[1] <=32'h3F0A5142;
	Rot_Kappa_Cir[2] <=32'h3F0A5142;
	Rot_Kappa_Cir[3] <=32'h3F0A5142;
	Rot_Kappa_Cir[4] <=32'h3F0A5142;
	Rot_Kappa_Cir[5] <=32'h3F0A5142;
	Rot_Kappa_Cir[6] <=32'h3F0A5142;
	Rot_Kappa_Cir[7] <=32'h3F0A5142;
	Rot_Kappa_Cir[8] <=32'h3F0A5142;
	Rot_Kappa_Cir[9] <=32'h3F0A5142;
	Rot_Kappa_Cir[10] <=32'h3F0A5142;
	Rot_Kappa_Cir[11] <=32'h3F0A5142;
	Rot_Kappa_Cir[12] <=32'h3F0A5142;
	Rot_Kappa_Cir[13] <=32'h3F0A5142;
	Rot_Kappa_Cir[14] <=32'h3F0A5142;
	Rot_Kappa_Cir[15] <=32'h3F0A5142;
	Rot_Kappa_Cir[16] <=32'h3F60A941;
	Rot_Kappa_Cir[17] <=32'h3F5CB779;
	Rot_Kappa_Cir[18] <=32'h3F588E83;
	Rot_Kappa_Cir[19] <=32'h3F542F6B;
	Rot_Kappa_Cir[20] <=32'h3F4F9B49;
	Rot_Kappa_Cir[21] <=32'h3F4AD340;
	Rot_Kappa_Cir[22] <=32'h3F45D884;
	Rot_Kappa_Cir[23] <=32'h3F40AC53;
	Rot_Kappa_Cir[24] <=32'h3F3B4FF7;
	Rot_Kappa_Cir[25] <=32'h3F35C4C9;
	Rot_Kappa_Cir[26] <=32'h3F300C2A;
	Rot_Kappa_Cir[27] <=32'h3F2A278A;
	Rot_Kappa_Cir[28] <=32'h3F241860;
	Rot_Kappa_Cir[29] <=32'h3F1DE031;
	Rot_Kappa_Cir[30] <=32'h3F17808B;
	Rot_Kappa_Cir[31] <=32'h3F10FB05;
	Rot_Kappa_Cir[32] <=32'h3F780AA6;
	Rot_Kappa_Cir[33] <=32'h3F770591;
	Rot_Kappa_Cir[34] <=32'h3F75F10C;
	Rot_Kappa_Cir[35] <=32'h3F74CD27;
	Rot_Kappa_Cir[36] <=32'h3F7399F6;
	Rot_Kappa_Cir[37] <=32'h3F72578C;
	Rot_Kappa_Cir[38] <=32'h3F7105FB;
	Rot_Kappa_Cir[39] <=32'h3F6FA55B;
	Rot_Kappa_Cir[40] <=32'h3F6E35C1;
	Rot_Kappa_Cir[41] <=32'h3F6CB743;
	Rot_Kappa_Cir[42] <=32'h3F6B29F9;
	Rot_Kappa_Cir[43] <=32'h3F698DFE;
	Rot_Kappa_Cir[44] <=32'h3F67E369;
	Rot_Kappa_Cir[45] <=32'h3F662A56;
	Rot_Kappa_Cir[46] <=32'h3F6462E1;
	Rot_Kappa_Cir[47] <=32'h3F628D26;
	Rot_Kappa_Cir[48] <=32'h3F7E00AC;
	Rot_Kappa_Cir[49] <=32'h3F7DBEDB;
	Rot_Kappa_Cir[50] <=32'h3F7D7912;
	Rot_Kappa_Cir[51] <=32'h3F7D2F54;
	Rot_Kappa_Cir[52] <=32'h3F7CE1A2;
	Rot_Kappa_Cir[53] <=32'h3F7C8FFB;
	Rot_Kappa_Cir[54] <=32'h3F7C3A63;
	Rot_Kappa_Cir[55] <=32'h3F7BE0D9;
	Rot_Kappa_Cir[56] <=32'h3F7B8360;
	Rot_Kappa_Cir[57] <=32'h3F7B21F9;
	Rot_Kappa_Cir[58] <=32'h3F7ABCA6;
	Rot_Kappa_Cir[59] <=32'h3F7A5367;
	Rot_Kappa_Cir[60] <=32'h3F79E63F;
	Rot_Kappa_Cir[61] <=32'h3F797530;
	Rot_Kappa_Cir[62] <=32'h3F79003B;
	Rot_Kappa_Cir[63] <=32'h3F788761;
	Rot_Kappa_Cir[64] <=32'h3F7F800C;
	Rot_Kappa_Cir[65] <=32'h3F7F6F8F;
	Rot_Kappa_Cir[66] <=32'h3F7F5E12;
	Rot_Kappa_Cir[67] <=32'h3F7F4B96;
	Rot_Kappa_Cir[68] <=32'h3F7F381B;
	Rot_Kappa_Cir[69] <=32'h3F7F23A1;
	Rot_Kappa_Cir[70] <=32'h3F7F0E27;
	Rot_Kappa_Cir[71] <=32'h3F7EF7AF;
	Rot_Kappa_Cir[72] <=32'h3F7EE037;
	Rot_Kappa_Cir[73] <=32'h3F7EC7C1;
	Rot_Kappa_Cir[74] <=32'h3F7EAE4C;
	Rot_Kappa_Cir[75] <=32'h3F7E93D8;
	Rot_Kappa_Cir[76] <=32'h3F7E7865;
	Rot_Kappa_Cir[77] <=32'h3F7E5BF4;
	Rot_Kappa_Cir[78] <=32'h3F7E3E85;
	Rot_Kappa_Cir[79] <=32'h3F7E2017;
	Rot_Kappa_Cir[80] <=32'h3F7FE002;
	Rot_Kappa_Cir[81] <=32'h3F7FDBE2;
	Rot_Kappa_Cir[82] <=32'h3F7FD782;
	Rot_Kappa_Cir[83] <=32'h3F7FD2E3;
	Rot_Kappa_Cir[84] <=32'h3F7FCE03;
	Rot_Kappa_Cir[85] <=32'h3F7FC8E3;
	Rot_Kappa_Cir[86] <=32'h3F7FC384;
	Rot_Kappa_Cir[87] <=32'h3F7FBDE4;
	Rot_Kappa_Cir[88] <=32'h3F7FB805;
	Rot_Kappa_Cir[89] <=32'h3F7FB1E5;
	Rot_Kappa_Cir[90] <=32'h3F7FAB86;
	Rot_Kappa_Cir[91] <=32'h3F7FA4E7;
	Rot_Kappa_Cir[92] <=32'h3F7F9E07;
	Rot_Kappa_Cir[93] <=32'h3F7F96E8;
	Rot_Kappa_Cir[94] <=32'h3F7F8F89;
	Rot_Kappa_Cir[95] <=32'h3F7F87EB;
	Rot_Kappa_Cir[96] <=32'h3F7FF801;
	Rot_Kappa_Cir[97] <=32'h3F7FF6F9;
	Rot_Kappa_Cir[98] <=32'h3F7FF5E1;
	Rot_Kappa_Cir[99] <=32'h3F7FF4B9;
	Rot_Kappa_Cir[100] <=32'h3F7FF381;
	Rot_Kappa_Cir[101] <=32'h3F7FF239;
	Rot_Kappa_Cir[102] <=32'h3F7FF0E1;
	Rot_Kappa_Cir[103] <=32'h3F7FEF79;
	Rot_Kappa_Cir[104] <=32'h3F7FEE01;
	Rot_Kappa_Cir[105] <=32'h3F7FEC79;
	Rot_Kappa_Cir[106] <=32'h3F7FEAE1;
	Rot_Kappa_Cir[107] <=32'h3F7FE93A;
	Rot_Kappa_Cir[108] <=32'h3F7FE782;
	Rot_Kappa_Cir[109] <=32'h3F7FE5BA;
	Rot_Kappa_Cir[110] <=32'h3F7FE3E2;
	Rot_Kappa_Cir[111] <=32'h3F7FE1FA;
	Rot_Kappa_Cir[112] <=32'h3F7FFE01;
	Rot_Kappa_Cir[113] <=32'h3F7FFDBF;
	Rot_Kappa_Cir[114] <=32'h3F7FFD79;
	Rot_Kappa_Cir[115] <=32'h3F7FFD2F;
	Rot_Kappa_Cir[116] <=32'h3F7FFCE1;
	Rot_Kappa_Cir[117] <=32'h3F7FFC8F;
	Rot_Kappa_Cir[118] <=32'h3F7FFC39;
	Rot_Kappa_Cir[119] <=32'h3F7FFBDF;
	Rot_Kappa_Cir[120] <=32'h3F7FFB81;
	Rot_Kappa_Cir[121] <=32'h3F7FFB1F;
	Rot_Kappa_Cir[122] <=32'h3F7FFAB9;
	Rot_Kappa_Cir[123] <=32'h3F7FFA4F;
	Rot_Kappa_Cir[124] <=32'h3F7FF9E1;
	Rot_Kappa_Cir[125] <=32'h3F7FF96F;
	Rot_Kappa_Cir[126] <=32'h3F7FF8F9;
	Rot_Kappa_Cir[127] <=32'h3F7FF87F;
	Rot_Kappa_Cir[128] <=32'h3F7FFF81;
	Rot_Kappa_Cir[129] <=32'h3F7FFF71;
	Rot_Kappa_Cir[130] <=32'h3F7FFF5F;
	Rot_Kappa_Cir[131] <=32'h3F7FFF4D;
	Rot_Kappa_Cir[132] <=32'h3F7FFF39;
	Rot_Kappa_Cir[133] <=32'h3F7FFF25;
	Rot_Kappa_Cir[134] <=32'h3F7FFF0F;
	Rot_Kappa_Cir[135] <=32'h3F7FFEF9;
	Rot_Kappa_Cir[136] <=32'h3F7FFEE1;
	Rot_Kappa_Cir[137] <=32'h3F7FFEC9;
	Rot_Kappa_Cir[138] <=32'h3F7FFEAF;
	Rot_Kappa_Cir[139] <=32'h3F7FFE95;
	Rot_Kappa_Cir[140] <=32'h3F7FFE79;
	Rot_Kappa_Cir[141] <=32'h3F7FFE5D;
	Rot_Kappa_Cir[142] <=32'h3F7FFE3F;
	Rot_Kappa_Cir[143] <=32'h3F7FFE21;
	Rot_Kappa_Cir[144] <=32'h3F7FFFE1;
	Rot_Kappa_Cir[145] <=32'h3F7FFFDD;
	Rot_Kappa_Cir[146] <=32'h3F7FFFD9;
	Rot_Kappa_Cir[147] <=32'h3F7FFFD4;
	Rot_Kappa_Cir[148] <=32'h3F7FFFCF;
	Rot_Kappa_Cir[149] <=32'h3F7FFFCA;
	Rot_Kappa_Cir[150] <=32'h3F7FFFC5;
	Rot_Kappa_Cir[151] <=32'h3F7FFFBF;
	Rot_Kappa_Cir[152] <=32'h3F7FFFB9;
	Rot_Kappa_Cir[153] <=32'h3F7FFFB3;
	Rot_Kappa_Cir[154] <=32'h3F7FFFAD;
	Rot_Kappa_Cir[155] <=32'h3F7FFFA6;
	Rot_Kappa_Cir[156] <=32'h3F7FFF9F;
	Rot_Kappa_Cir[157] <=32'h3F7FFF98;
	Rot_Kappa_Cir[158] <=32'h3F7FFF91;
	Rot_Kappa_Cir[159] <=32'h3F7FFF89;
	Rot_Kappa_Cir[160] <=32'h3F7FFFF9;
	Rot_Kappa_Cir[161] <=32'h3F7FFFF8;
	Rot_Kappa_Cir[162] <=32'h3F7FFFF7;
	Rot_Kappa_Cir[163] <=32'h3F7FFFF6;
	Rot_Kappa_Cir[164] <=32'h3F7FFFF5;
	Rot_Kappa_Cir[165] <=32'h3F7FFFF3;
	Rot_Kappa_Cir[166] <=32'h3F7FFFF2;
	Rot_Kappa_Cir[167] <=32'h3F7FFFF1;
	Rot_Kappa_Cir[168] <=32'h3F7FFFEF;
	Rot_Kappa_Cir[169] <=32'h3F7FFFEE;
	Rot_Kappa_Cir[170] <=32'h3F7FFFEC;
	Rot_Kappa_Cir[171] <=32'h3F7FFFEA;
	Rot_Kappa_Cir[172] <=32'h3F7FFFE9;
	Rot_Kappa_Cir[173] <=32'h3F7FFFE7;
	Rot_Kappa_Cir[174] <=32'h3F7FFFE5;
	Rot_Kappa_Cir[175] <=32'h3F7FFFE3;
	Rot_Kappa_Cir[176] <=32'h3F7FFFFF;
	Rot_Kappa_Cir[177] <=32'h3F7FFFFF;
	Rot_Kappa_Cir[178] <=32'h3F7FFFFF;
	Rot_Kappa_Cir[179] <=32'h3F7FFFFE;
	Rot_Kappa_Cir[180] <=32'h3F7FFFFE;
	Rot_Kappa_Cir[181] <=32'h3F7FFFFE;
	Rot_Kappa_Cir[182] <=32'h3F7FFFFD;
	Rot_Kappa_Cir[183] <=32'h3F7FFFFD;
	Rot_Kappa_Cir[184] <=32'h3F7FFFFD;
	Rot_Kappa_Cir[185] <=32'h3F7FFFFC;
	Rot_Kappa_Cir[186] <=32'h3F7FFFFC;
	Rot_Kappa_Cir[187] <=32'h3F7FFFFB;
	Rot_Kappa_Cir[188] <=32'h3F7FFFFB;
	Rot_Kappa_Cir[189] <=32'h3F7FFFFB;
	Rot_Kappa_Cir[190] <=32'h3F7FFFFA;
	Rot_Kappa_Cir[191] <=32'h3F7FFFFA;
	Rot_Kappa_Cir[192] <=32'h3F800000;
	Rot_Kappa_Cir[193] <=32'h3F800000;
	Rot_Kappa_Cir[194] <=32'h3F800000;
	Rot_Kappa_Cir[195] <=32'h3F800000;
	Rot_Kappa_Cir[196] <=32'h3F800000;
	Rot_Kappa_Cir[197] <=32'h3F800000;
	Rot_Kappa_Cir[198] <=32'h3F800000;
	Rot_Kappa_Cir[199] <=32'h3F800000;
	Rot_Kappa_Cir[200] <=32'h3F800000;
	Rot_Kappa_Cir[201] <=32'h3F800000;
	Rot_Kappa_Cir[202] <=32'h3F800000;
	Rot_Kappa_Cir[203] <=32'h3F800000;
	Rot_Kappa_Cir[204] <=32'h3F800000;
	Rot_Kappa_Cir[205] <=32'h3F800000;
	Rot_Kappa_Cir[206] <=32'h3F7FFFFF;
	Rot_Kappa_Cir[207] <=32'h3F7FFFFF;
	Rot_Kappa_Cir[208] <=32'h3F800000;
	Rot_Kappa_Cir[209] <=32'h3F800000;
	Rot_Kappa_Cir[210] <=32'h3F800000;
	Rot_Kappa_Cir[211] <=32'h3F800000;
	Rot_Kappa_Cir[212] <=32'h3F800000;
	Rot_Kappa_Cir[213] <=32'h3F800000;
	Rot_Kappa_Cir[214] <=32'h3F800000;
	Rot_Kappa_Cir[215] <=32'h3F800000;
	Rot_Kappa_Cir[216] <=32'h3F800000;
	Rot_Kappa_Cir[217] <=32'h3F800000;
	Rot_Kappa_Cir[218] <=32'h3F800000;
	Rot_Kappa_Cir[219] <=32'h3F800000;
	Rot_Kappa_Cir[220] <=32'h3F800000;
	Rot_Kappa_Cir[221] <=32'h3F800000;
	Rot_Kappa_Cir[222] <=32'h3F800000;
	Rot_Kappa_Cir[223] <=32'h3F800000;
	Rot_Kappa_Cir[224] <=32'h3F800000;
	Rot_Kappa_Cir[225] <=32'h3F800000;
	Rot_Kappa_Cir[226] <=32'h3F800000;
	Rot_Kappa_Cir[227] <=32'h3F800000;
	Rot_Kappa_Cir[228] <=32'h3F800000;
	Rot_Kappa_Cir[229] <=32'h3F800000;
	Rot_Kappa_Cir[230] <=32'h3F800000;
	Rot_Kappa_Cir[231] <=32'h3F800000;
	Rot_Kappa_Cir[232] <=32'h3F800000;
	Rot_Kappa_Cir[233] <=32'h3F800000;
	Rot_Kappa_Cir[234] <=32'h3F800000;
	Rot_Kappa_Cir[235] <=32'h3F800000;
	Rot_Kappa_Cir[236] <=32'h3F800000;
	Rot_Kappa_Cir[237] <=32'h3F800000;
	Rot_Kappa_Cir[238] <=32'h3F800000;
	Rot_Kappa_Cir[239] <=32'h3F800000;
	Rot_Kappa_Cir[240] <=32'h3F800000;
	Rot_Kappa_Cir[241] <=32'h3F800000;
	Rot_Kappa_Cir[242] <=32'h3F800000;
	Rot_Kappa_Cir[243] <=32'h3F800000;
	Rot_Kappa_Cir[244] <=32'h3F800000;
	Rot_Kappa_Cir[245] <=32'h3F800000;
	Rot_Kappa_Cir[246] <=32'h3F800000;
	Rot_Kappa_Cir[247] <=32'h3F800000;
	Rot_Kappa_Cir[248] <=32'h3F800000;
	Rot_Kappa_Cir[249] <=32'h3F800000;
	Rot_Kappa_Cir[250] <=32'h3F800000;
	Rot_Kappa_Cir[251] <=32'h3F800000;
	Rot_Kappa_Cir[252] <=32'h3F800000;
	Rot_Kappa_Cir[253] <=32'h3F800000;
	Rot_Kappa_Cir[254] <=32'h3F800000;
	Rot_Kappa_Cir[255] <=32'h3F800000;
	
	//Rotation Kappa Hyperbolic
	Rot_Kappa_Hyper[0] <=32'h3FC583AB;
	Rot_Kappa_Hyper[1] <=32'h3FCF4ED6;
	Rot_Kappa_Hyper[2] <=32'h3FD9E961;
	Rot_Kappa_Hyper[3] <=32'h3FE55DE8;
	Rot_Kappa_Hyper[4] <=32'h3FF1B7E0;
	Rot_Kappa_Hyper[5] <=32'h3FFF03A4;
	Rot_Kappa_Hyper[6] <=32'h4006A740;
	Rot_Kappa_Hyper[7] <=32'h400E5361;
	Rot_Kappa_Hyper[8] <=32'h40168DE1;
	Rot_Kappa_Hyper[9] <=32'h401F5EFB;
	Rot_Kappa_Hyper[10] <=32'h4028CF82;
	Rot_Kappa_Hyper[11] <=32'h4032E8E7;
	Rot_Kappa_Hyper[12] <=32'h403DB543;
	Rot_Kappa_Hyper[13] <=32'h40493F64;
	Rot_Kappa_Hyper[14] <=32'h405592D5;
	Rot_Kappa_Hyper[15] <=32'h4062BBEB;
	Rot_Kappa_Hyper[16] <=32'h3F90560D;
	Rot_Kappa_Hyper[17] <=32'h3F927DC8;
	Rot_Kappa_Hyper[18] <=32'h3F94CA23;
	Rot_Kappa_Hyper[19] <=32'h3F973BB2;
	Rot_Kappa_Hyper[20] <=32'h3F99D311;
	Rot_Kappa_Hyper[21] <=32'h3F9C90E5;
	Rot_Kappa_Hyper[22] <=32'h3F9F75DE;
	Rot_Kappa_Hyper[23] <=32'h3FA282B6;
	Rot_Kappa_Hyper[24] <=32'h3FA5B82F;
	Rot_Kappa_Hyper[25] <=32'h3FA91717;
	Rot_Kappa_Hyper[26] <=32'h3FACA045;
	Rot_Kappa_Hyper[27] <=32'h3FB0549D;
	Rot_Kappa_Hyper[28] <=32'h3FB4350B;
	Rot_Kappa_Hyper[29] <=32'h3FB84286;
	Rot_Kappa_Hyper[30] <=32'h3FBC7E14;
	Rot_Kappa_Hyper[31] <=32'h3FC0E8C2;
	Rot_Kappa_Hyper[32] <=32'h3F840559;
	Rot_Kappa_Hyper[33] <=32'h3F848AD0;
	Rot_Kappa_Hyper[34] <=32'h3F851891;
	Rot_Kappa_Hyper[35] <=32'h3F85AEA3;
	Rot_Kappa_Hyper[36] <=32'h3F864D11;
	Rot_Kappa_Hyper[37] <=32'h3F86F3E3;
	Rot_Kappa_Hyper[38] <=32'h3F87A324;
	Rot_Kappa_Hyper[39] <=32'h3F885AE0;
	Rot_Kappa_Hyper[40] <=32'h3F891B21;
	Rot_Kappa_Hyper[41] <=32'h3F89E3F4;
	Rot_Kappa_Hyper[42] <=32'h3F8AB565;
	Rot_Kappa_Hyper[43] <=32'h3F8B8F82;
	Rot_Kappa_Hyper[44] <=32'h3F8C7258;
	Rot_Kappa_Hyper[45] <=32'h3F8D5DF5;
	Rot_Kappa_Hyper[46] <=32'h3F8E5267;
	Rot_Kappa_Hyper[47] <=32'h3F8F4FBF;
	Rot_Kappa_Hyper[48] <=32'h3F810056;
	Rot_Kappa_Hyper[49] <=32'h3F81216D;
	Rot_Kappa_Hyper[50] <=32'h3F814489;
	Rot_Kappa_Hyper[51] <=32'h3F8169AA;
	Rot_Kappa_Hyper[52] <=32'h3F8190D1;
	Rot_Kappa_Hyper[53] <=32'h3F81B9FE;
	Rot_Kappa_Hyper[54] <=32'h3F81E532;
	Rot_Kappa_Hyper[55] <=32'h3F82126D;
	Rot_Kappa_Hyper[56] <=32'h3F8241B1;
	Rot_Kappa_Hyper[57] <=32'h3F8272FE;
	Rot_Kappa_Hyper[58] <=32'h3F82A654;
	Rot_Kappa_Hyper[59] <=32'h3F82DBB5;
	Rot_Kappa_Hyper[60] <=32'h3F831322;
	Rot_Kappa_Hyper[61] <=32'h3F834C9B;
	Rot_Kappa_Hyper[62] <=32'h3F838821;
	Rot_Kappa_Hyper[63] <=32'h3F83C5B5;
	Rot_Kappa_Hyper[64] <=32'h3F804006;
	Rot_Kappa_Hyper[65] <=32'h3F804847;
	Rot_Kappa_Hyper[66] <=32'h3F805109;
	Rot_Kappa_Hyper[67] <=32'h3F805A4B;
	Rot_Kappa_Hyper[68] <=32'h3F80640D;
	Rot_Kappa_Hyper[69] <=32'h3F806E50;
	Rot_Kappa_Hyper[70] <=32'h3F807913;
	Rot_Kappa_Hyper[71] <=32'h3F808457;
	Rot_Kappa_Hyper[72] <=32'h3F80901B;
	Rot_Kappa_Hyper[73] <=32'h3F809C60;
	Rot_Kappa_Hyper[74] <=32'h3F80A926;
	Rot_Kappa_Hyper[75] <=32'h3F80B66C;
	Rot_Kappa_Hyper[76] <=32'h3F80C432;
	Rot_Kappa_Hyper[77] <=32'h3F80D27A;
	Rot_Kappa_Hyper[78] <=32'h3F80E142;
	Rot_Kappa_Hyper[79] <=32'h3F80F08C;
	Rot_Kappa_Hyper[80] <=32'h3F801001;
	Rot_Kappa_Hyper[81] <=32'h3F801211;
	Rot_Kappa_Hyper[82] <=32'h3F801441;
	Rot_Kappa_Hyper[83] <=32'h3F801691;
	Rot_Kappa_Hyper[84] <=32'h3F801901;
	Rot_Kappa_Hyper[85] <=32'h3F801B91;
	Rot_Kappa_Hyper[86] <=32'h3F801E42;
	Rot_Kappa_Hyper[87] <=32'h3F802112;
	Rot_Kappa_Hyper[88] <=32'h3F802402;
	Rot_Kappa_Hyper[89] <=32'h3F802712;
	Rot_Kappa_Hyper[90] <=32'h3F802A43;
	Rot_Kappa_Hyper[91] <=32'h3F802D93;
	Rot_Kappa_Hyper[92] <=32'h3F803103;
	Rot_Kappa_Hyper[93] <=32'h3F803494;
	Rot_Kappa_Hyper[94] <=32'h3F803844;
	Rot_Kappa_Hyper[95] <=32'h3F803C15;
	Rot_Kappa_Hyper[96] <=32'h3F800400;
	Rot_Kappa_Hyper[97] <=32'h3F800484;
	Rot_Kappa_Hyper[98] <=32'h3F800510;
	Rot_Kappa_Hyper[99] <=32'h3F8005A4;
	Rot_Kappa_Hyper[100] <=32'h3F800640;
	Rot_Kappa_Hyper[101] <=32'h3F8006E4;
	Rot_Kappa_Hyper[102] <=32'h3F800790;
	Rot_Kappa_Hyper[103] <=32'h3F800844;
	Rot_Kappa_Hyper[104] <=32'h3F800900;
	Rot_Kappa_Hyper[105] <=32'h3F8009C4;
	Rot_Kappa_Hyper[106] <=32'h3F800A90;
	Rot_Kappa_Hyper[107] <=32'h3F800B65;
	Rot_Kappa_Hyper[108] <=32'h3F800C41;
	Rot_Kappa_Hyper[109] <=32'h3F800D25;
	Rot_Kappa_Hyper[110] <=32'h3F800E11;
	Rot_Kappa_Hyper[111] <=32'h3F800F05;
	Rot_Kappa_Hyper[112] <=32'h3F800100;
	Rot_Kappa_Hyper[113] <=32'h3F800121;
	Rot_Kappa_Hyper[114] <=32'h3F800144;
	Rot_Kappa_Hyper[115] <=32'h3F800169;
	Rot_Kappa_Hyper[116] <=32'h3F800190;
	Rot_Kappa_Hyper[117] <=32'h3F8001B9;
	Rot_Kappa_Hyper[118] <=32'h3F8001E4;
	Rot_Kappa_Hyper[119] <=32'h3F800211;
	Rot_Kappa_Hyper[120] <=32'h3F800240;
	Rot_Kappa_Hyper[121] <=32'h3F800271;
	Rot_Kappa_Hyper[122] <=32'h3F8002A4;
	Rot_Kappa_Hyper[123] <=32'h3F8002D9;
	Rot_Kappa_Hyper[124] <=32'h3F800310;
	Rot_Kappa_Hyper[125] <=32'h3F800349;
	Rot_Kappa_Hyper[126] <=32'h3F800384;
	Rot_Kappa_Hyper[127] <=32'h3F8003C1;
	Rot_Kappa_Hyper[128] <=32'h3F800040;
	Rot_Kappa_Hyper[129] <=32'h3F800049;
	Rot_Kappa_Hyper[130] <=32'h3F800051;
	Rot_Kappa_Hyper[131] <=32'h3F80005B;
	Rot_Kappa_Hyper[132] <=32'h3F800064;
	Rot_Kappa_Hyper[133] <=32'h3F80006F;
	Rot_Kappa_Hyper[134] <=32'h3F800079;
	Rot_Kappa_Hyper[135] <=32'h3F800085;
	Rot_Kappa_Hyper[136] <=32'h3F800090;
	Rot_Kappa_Hyper[137] <=32'h3F80009D;
	Rot_Kappa_Hyper[138] <=32'h3F8000A9;
	Rot_Kappa_Hyper[139] <=32'h3F8000B7;
	Rot_Kappa_Hyper[140] <=32'h3F8000C4;
	Rot_Kappa_Hyper[141] <=32'h3F8000D3;
	Rot_Kappa_Hyper[142] <=32'h3F8000E1;
	Rot_Kappa_Hyper[143] <=32'h3F8000F1;
	Rot_Kappa_Hyper[144] <=32'h3F800010;
	Rot_Kappa_Hyper[145] <=32'h3F800012;
	Rot_Kappa_Hyper[146] <=32'h3F800015;
	Rot_Kappa_Hyper[147] <=32'h3F800017;
	Rot_Kappa_Hyper[148] <=32'h3F800019;
	Rot_Kappa_Hyper[149] <=32'h3F80001C;
	Rot_Kappa_Hyper[150] <=32'h3F80001F;
	Rot_Kappa_Hyper[151] <=32'h3F800021;
	Rot_Kappa_Hyper[152] <=32'h3F800024;
	Rot_Kappa_Hyper[153] <=32'h3F800027;
	Rot_Kappa_Hyper[154] <=32'h3F80002B;
	Rot_Kappa_Hyper[155] <=32'h3F80002E;
	Rot_Kappa_Hyper[156] <=32'h3F800031;
	Rot_Kappa_Hyper[157] <=32'h3F800035;
	Rot_Kappa_Hyper[158] <=32'h3F800039;
	Rot_Kappa_Hyper[159] <=32'h3F80003C;
	Rot_Kappa_Hyper[160] <=32'h3F800004;
	Rot_Kappa_Hyper[161] <=32'h3F800005;
	Rot_Kappa_Hyper[162] <=32'h3F800005;
	Rot_Kappa_Hyper[163] <=32'h3F800006;
	Rot_Kappa_Hyper[164] <=32'h3F800007;
	Rot_Kappa_Hyper[165] <=32'h3F800007;
	Rot_Kappa_Hyper[166] <=32'h3F800008;
	Rot_Kappa_Hyper[167] <=32'h3F800009;
	Rot_Kappa_Hyper[168] <=32'h3F800009;
	Rot_Kappa_Hyper[169] <=32'h3F80000A;
	Rot_Kappa_Hyper[170] <=32'h3F80000B;
	Rot_Kappa_Hyper[171] <=32'h3F80000C;
	Rot_Kappa_Hyper[172] <=32'h3F80000D;
	Rot_Kappa_Hyper[173] <=32'h3F80000D;
	Rot_Kappa_Hyper[174] <=32'h3F80000E;
	Rot_Kappa_Hyper[175] <=32'h3F80000F;
	Rot_Kappa_Hyper[176] <=32'h3F800001;
	Rot_Kappa_Hyper[177] <=32'h3F800001;
	Rot_Kappa_Hyper[178] <=32'h3F800002;
	Rot_Kappa_Hyper[179] <=32'h3F800002;
	Rot_Kappa_Hyper[180] <=32'h3F800002;
	Rot_Kappa_Hyper[181] <=32'h3F800002;
	Rot_Kappa_Hyper[182] <=32'h3F800002;
	Rot_Kappa_Hyper[183] <=32'h3F800002;
	Rot_Kappa_Hyper[184] <=32'h3F800003;
	Rot_Kappa_Hyper[185] <=32'h3F800003;
	Rot_Kappa_Hyper[186] <=32'h3F800003;
	Rot_Kappa_Hyper[187] <=32'h3F800003;
	Rot_Kappa_Hyper[188] <=32'h3F800003;
	Rot_Kappa_Hyper[189] <=32'h3F800004;
	Rot_Kappa_Hyper[190] <=32'h3F800004;
	Rot_Kappa_Hyper[191] <=32'h3F800004;
	Rot_Kappa_Hyper[192] <=32'h3F800001;
	Rot_Kappa_Hyper[193] <=32'h3F800001;
	Rot_Kappa_Hyper[194] <=32'h3F800001;
	Rot_Kappa_Hyper[195] <=32'h3F800001;
	Rot_Kappa_Hyper[196] <=32'h3F800001;
	Rot_Kappa_Hyper[197] <=32'h3F800001;
	Rot_Kappa_Hyper[198] <=32'h3F800001;
	Rot_Kappa_Hyper[199] <=32'h3F800001;
	Rot_Kappa_Hyper[200] <=32'h3F800001;
	Rot_Kappa_Hyper[201] <=32'h3F800001;
	Rot_Kappa_Hyper[202] <=32'h3F800001;
	Rot_Kappa_Hyper[203] <=32'h3F800001;
	Rot_Kappa_Hyper[204] <=32'h3F800001;
	Rot_Kappa_Hyper[205] <=32'h3F800001;
	Rot_Kappa_Hyper[206] <=32'h3F800001;
	Rot_Kappa_Hyper[207] <=32'h3F800001;
	Rot_Kappa_Hyper[208] <=32'h3F800000;
	Rot_Kappa_Hyper[209] <=32'h3F800000;
	Rot_Kappa_Hyper[210] <=32'h3F800000;
	Rot_Kappa_Hyper[211] <=32'h3F800000;
	Rot_Kappa_Hyper[212] <=32'h3F800000;
	Rot_Kappa_Hyper[213] <=32'h3F800000;
	Rot_Kappa_Hyper[214] <=32'h3F800000;
	Rot_Kappa_Hyper[215] <=32'h3F800000;
	Rot_Kappa_Hyper[216] <=32'h3F800000;
	Rot_Kappa_Hyper[217] <=32'h3F800000;
	Rot_Kappa_Hyper[218] <=32'h3F800001;
	Rot_Kappa_Hyper[219] <=32'h3F800001;
	Rot_Kappa_Hyper[220] <=32'h3F800001;
	Rot_Kappa_Hyper[221] <=32'h3F800001;
	Rot_Kappa_Hyper[222] <=32'h3F800001;
	Rot_Kappa_Hyper[223] <=32'h3F800001;
	Rot_Kappa_Hyper[224] <=32'h3F800000;
	Rot_Kappa_Hyper[225] <=32'h3F800000;
	Rot_Kappa_Hyper[226] <=32'h3F800000;
	Rot_Kappa_Hyper[227] <=32'h3F800000;
	Rot_Kappa_Hyper[228] <=32'h3F800000;
	Rot_Kappa_Hyper[229] <=32'h3F800000;
	Rot_Kappa_Hyper[230] <=32'h3F800000;
	Rot_Kappa_Hyper[231] <=32'h3F800000;
	Rot_Kappa_Hyper[232] <=32'h3F800000;
	Rot_Kappa_Hyper[233] <=32'h3F800000;
	Rot_Kappa_Hyper[234] <=32'h3F800000;
	Rot_Kappa_Hyper[235] <=32'h3F800000;
	Rot_Kappa_Hyper[236] <=32'h3F800000;
	Rot_Kappa_Hyper[237] <=32'h3F800000;
	Rot_Kappa_Hyper[238] <=32'h3F800000;
	Rot_Kappa_Hyper[239] <=32'h3F800000;
	Rot_Kappa_Hyper[240] <=32'h3F800000;
	Rot_Kappa_Hyper[241] <=32'h3F800000;
	Rot_Kappa_Hyper[242] <=32'h3F800000;
	Rot_Kappa_Hyper[243] <=32'h3F800000;
	Rot_Kappa_Hyper[244] <=32'h3F800000;
	Rot_Kappa_Hyper[245] <=32'h3F800000;
	Rot_Kappa_Hyper[246] <=32'h3F800000;
	Rot_Kappa_Hyper[247] <=32'h3F800000;
	Rot_Kappa_Hyper[248] <=32'h3F800000;
	Rot_Kappa_Hyper[249] <=32'h3F800000;
	Rot_Kappa_Hyper[250] <=32'h3F800000;
	Rot_Kappa_Hyper[251] <=32'h3F800000;
	Rot_Kappa_Hyper[252] <=32'h3F800000;
	Rot_Kappa_Hyper[253] <=32'h3F800000;
	Rot_Kappa_Hyper[254] <=32'h3F800000;
	Rot_Kappa_Hyper[255] <=32'h3F800000;

	// Delta vectoring
	Vec_Delta[0] <=32'h3F4CCCDE;
	Vec_Delta[1] <=32'h3F2AAABC;
	Vec_Delta[2] <=32'h3F124936;
	Vec_Delta[3] <=32'h3F000011;
	Vec_Delta[4] <=32'h3F800009;
	Vec_Delta[5] <=32'h3F555567;
	Vec_Delta[6] <=32'h3F36DB7F;
	Vec_Delta[7] <=32'h3F200011;
	Vec_Delta[8] <=32'h3F9999A2;
	Vec_Delta[9] <=32'h3F800009;
	Vec_Delta[10] <=32'h3F5B6DC8;
	Vec_Delta[11] <=32'h3F400011;
	Vec_Delta[12] <=32'h3FB3333C;
	Vec_Delta[13] <=32'h3F95555E;
	Vec_Delta[14] <=32'h3F800008;
	Vec_Delta[15] <=32'h3F600011;
	Vec_Delta[16] <=32'h3ECCCCEF;
	Vec_Delta[17] <=32'h3EAAAACD;
	Vec_Delta[18] <=32'h3E924946;
	Vec_Delta[19] <=32'h3E800022;
	Vec_Delta[20] <=32'h3F000011;
	Vec_Delta[21] <=32'h3ED55577;
	Vec_Delta[22] <=32'h3EB6DB90;
	Vec_Delta[23] <=32'h3EA00022;
	Vec_Delta[24] <=32'h3F1999AB;
	Vec_Delta[25] <=32'h3F000011;
	Vec_Delta[26] <=32'h3EDB6DD9;
	Vec_Delta[27] <=32'h3EC00022;
	Vec_Delta[28] <=32'h3F333345;
	Vec_Delta[29] <=32'h3F155566;
	Vec_Delta[30] <=32'h3F000011;
	Vec_Delta[31] <=32'h3EE00022;
	Vec_Delta[32] <=32'h3E4CCD11;
	Vec_Delta[33] <=32'h3E2AAAEE;
	Vec_Delta[34] <=32'h3E124968;
	Vec_Delta[35] <=32'h3E000043;
	Vec_Delta[36] <=32'h3E800022;
	Vec_Delta[37] <=32'h3E555599;
	Vec_Delta[38] <=32'h3E36DBB1;
	Vec_Delta[39] <=32'h3E200043;
	Vec_Delta[40] <=32'h3E9999BC;
	Vec_Delta[41] <=32'h3E800022;
	Vec_Delta[42] <=32'h3E5B6DFA;
	Vec_Delta[43] <=32'h3E400043;
	Vec_Delta[44] <=32'h3EB33355;
	Vec_Delta[45] <=32'h3E955577;
	Vec_Delta[46] <=32'h3E800022;
	Vec_Delta[47] <=32'h3E600043;
	Vec_Delta[48] <=32'h3DCCCD54;
	Vec_Delta[49] <=32'h3DAAAB31;
	Vec_Delta[50] <=32'h3D9249AB;
	Vec_Delta[51] <=32'h3D800086;
	Vec_Delta[52] <=32'h3E000043;
	Vec_Delta[53] <=32'h3DD555DC;
	Vec_Delta[54] <=32'h3DB6DBF4;
	Vec_Delta[55] <=32'h3DA00086;
	Vec_Delta[56] <=32'h3E1999DD;
	Vec_Delta[57] <=32'h3E000043;
	Vec_Delta[58] <=32'h3DDB6E3E;
	Vec_Delta[59] <=32'h3DC00086;
	Vec_Delta[60] <=32'h3E333377;
	Vec_Delta[61] <=32'h3E155599;
	Vec_Delta[62] <=32'h3E000043;
	Vec_Delta[63] <=32'h3DE00087;
	Vec_Delta[64] <=32'h3D4CCDDA;
	Vec_Delta[65] <=32'h3D2AABB7;
	Vec_Delta[66] <=32'h3D124A31;
	Vec_Delta[67] <=32'h3D00010C;
	Vec_Delta[68] <=32'h3D800087;
	Vec_Delta[69] <=32'h3D555662;
	Vec_Delta[70] <=32'h3D36DC7A;
	Vec_Delta[71] <=32'h3D20010D;
	Vec_Delta[72] <=32'h3D999A20;
	Vec_Delta[73] <=32'h3D800086;
	Vec_Delta[74] <=32'h3D5B6EC4;
	Vec_Delta[75] <=32'h3D40010D;
	Vec_Delta[76] <=32'h3DB333BA;
	Vec_Delta[77] <=32'h3D9555DC;
	Vec_Delta[78] <=32'h3D800086;
	Vec_Delta[79] <=32'h3D60010D;
	Vec_Delta[80] <=32'h3CCCCEE6;
	Vec_Delta[81] <=32'h3CAAACC4;
	Vec_Delta[82] <=32'h3C924B3E;
	Vec_Delta[83] <=32'h3C800219;
	Vec_Delta[84] <=32'h3D00010D;
	Vec_Delta[85] <=32'h3CD5576F;
	Vec_Delta[86] <=32'h3CB6DD87;
	Vec_Delta[87] <=32'h3CA00219;
	Vec_Delta[88] <=32'h3D199AA6;
	Vec_Delta[89] <=32'h3D00010D;
	Vec_Delta[90] <=32'h3CDB6FD0;
	Vec_Delta[91] <=32'h3CC00219;
	Vec_Delta[92] <=32'h3D333440;
	Vec_Delta[93] <=32'h3D155662;
	Vec_Delta[94] <=32'h3D00010D;
	Vec_Delta[95] <=32'h3CE00219;
	Vec_Delta[96] <=32'h3C4CD0FF;
	Vec_Delta[97] <=32'h3C2AAEDD;
	Vec_Delta[98] <=32'h3C124D56;
	Vec_Delta[99] <=32'h3C000432;
	Vec_Delta[100] <=32'h3C800219;
	Vec_Delta[101] <=32'h3C555988;
	Vec_Delta[102] <=32'h3C36DFA0;
	Vec_Delta[103] <=32'h3C200432;
	Vec_Delta[104] <=32'h3C999BB3;
	Vec_Delta[105] <=32'h3C800219;
	Vec_Delta[106] <=32'h3C5B71E9;
	Vec_Delta[107] <=32'h3C400432;
	Vec_Delta[108] <=32'h3CB3354D;
	Vec_Delta[109] <=32'h3C95576E;
	Vec_Delta[110] <=32'h3C800219;
	Vec_Delta[111] <=32'h3C600432;
	Vec_Delta[112] <=32'h3BCCD531;
	Vec_Delta[113] <=32'h3BAAB30F;
	Vec_Delta[114] <=32'h3B925188;
	Vec_Delta[115] <=32'h3B800863;
	Vec_Delta[116] <=32'h3C000432;
	Vec_Delta[117] <=32'h3BD55DB9;
	Vec_Delta[118] <=32'h3BB6E3D2;
	Vec_Delta[119] <=32'h3BA00864;
	Vec_Delta[120] <=32'h3C199DCC;
	Vec_Delta[121] <=32'h3C000432;
	Vec_Delta[122] <=32'h3BDB761B;
	Vec_Delta[123] <=32'h3BC00864;
	Vec_Delta[124] <=32'h3C333766;
	Vec_Delta[125] <=32'h3C155987;
	Vec_Delta[126] <=32'h3C000432;
	Vec_Delta[127] <=32'h3BE00864;
	Vec_Delta[128] <=32'h3B4CDD95;
	Vec_Delta[129] <=32'h3B2ABB72;
	Vec_Delta[130] <=32'h3B1259EC;
	Vec_Delta[131] <=32'h3B0010C7;
	Vec_Delta[132] <=32'h3B800864;
	Vec_Delta[133] <=32'h3B55661D;
	Vec_Delta[134] <=32'h3B36EC35;
	Vec_Delta[135] <=32'h3B2010C7;
	Vec_Delta[136] <=32'h3B99A1FE;
	Vec_Delta[137] <=32'h3B800864;
	Vec_Delta[138] <=32'h3B5B7E7E;
	Vec_Delta[139] <=32'h3B4010C7;
	Vec_Delta[140] <=32'h3BB33B97;
	Vec_Delta[141] <=32'h3B955DB9;
	Vec_Delta[142] <=32'h3B800864;
	Vec_Delta[143] <=32'h3B6010C7;
	Vec_Delta[144] <=32'h3ACCEE5C;
	Vec_Delta[145] <=32'h3AAACC39;
	Vec_Delta[146] <=32'h3A926AB3;
	Vec_Delta[147] <=32'h3A80218E;
	Vec_Delta[148] <=32'h3B0010C7;
	Vec_Delta[149] <=32'h3AD576E4;
	Vec_Delta[150] <=32'h3AB6FCFC;
	Vec_Delta[151] <=32'h3AA0218E;
	Vec_Delta[152] <=32'h3B19AA61;
	Vec_Delta[153] <=32'h3B0010C7;
	Vec_Delta[154] <=32'h3ADB8F45;
	Vec_Delta[155] <=32'h3AC0218E;
	Vec_Delta[156] <=32'h3B3343FB;
	Vec_Delta[157] <=32'h3B15661D;
	Vec_Delta[158] <=32'h3B0010C7;
	Vec_Delta[159] <=32'h3AE0218E;
	Vec_Delta[160] <=32'h3A4D0FE9;
	Vec_Delta[161] <=32'h3A2AEDC7;
	Vec_Delta[162] <=32'h3A128C41;
	Vec_Delta[163] <=32'h3A00431C;
	Vec_Delta[164] <=32'h3A80218E;
	Vec_Delta[165] <=32'h3A559872;
	Vec_Delta[166] <=32'h3A371E8A;
	Vec_Delta[167] <=32'h3A20431C;
	Vec_Delta[168] <=32'h3A99BB28;
	Vec_Delta[169] <=32'h3A80218E;
	Vec_Delta[170] <=32'h3A5BB0D3;
	Vec_Delta[171] <=32'h3A40431C;
	Vec_Delta[172] <=32'h3AB354C2;
	Vec_Delta[173] <=32'h3A9576E4;
	Vec_Delta[174] <=32'h3A80218E;
	Vec_Delta[175] <=32'h3A60431C;
	Vec_Delta[176] <=32'h39CD5305;
	Vec_Delta[177] <=32'h39AB30E3;
	Vec_Delta[178] <=32'h3992CF5C;
	Vec_Delta[179] <=32'h39808638;
	Vec_Delta[180] <=32'h3A00431C;
	Vec_Delta[181] <=32'h39D5DB8E;
	Vec_Delta[182] <=32'h39B761A6;
	Vec_Delta[183] <=32'h39A08638;
	Vec_Delta[184] <=32'h3A19DCB6;
	Vec_Delta[185] <=32'h3A00431C;
	Vec_Delta[186] <=32'h39DBF3EF;
	Vec_Delta[187] <=32'h39C08638;
	Vec_Delta[188] <=32'h3A337650;
	Vec_Delta[189] <=32'h3A159871;
	Vec_Delta[190] <=32'h3A00431C;
	Vec_Delta[191] <=32'h39E08638;
	Vec_Delta[192] <=32'h394DD93D;
	Vec_Delta[193] <=32'h392BB71B;
	Vec_Delta[194] <=32'h39135594;
	Vec_Delta[195] <=32'h39010C6F;
	Vec_Delta[196] <=32'h39808638;
	Vec_Delta[197] <=32'h395661C5;
	Vec_Delta[198] <=32'h3937E7DE;
	Vec_Delta[199] <=32'h39210C70;
	Vec_Delta[200] <=32'h399A1FD2;
	Vec_Delta[201] <=32'h39808638;
	Vec_Delta[202] <=32'h395C7A27;
	Vec_Delta[203] <=32'h39410C70;
	Vec_Delta[204] <=32'h39B3B96C;
	Vec_Delta[205] <=32'h3995DB8D;
	Vec_Delta[206] <=32'h39808638;
	Vec_Delta[207] <=32'h39610C70;
	Vec_Delta[208] <=32'h38CEE5AD;
	Vec_Delta[209] <=32'h38ACC38A;
	Vec_Delta[210] <=32'h38946204;
	Vec_Delta[211] <=32'h388218DF;
	Vec_Delta[212] <=32'h39010C70;
	Vec_Delta[213] <=32'h38D76E35;
	Vec_Delta[214] <=32'h38B8F44D;
	Vec_Delta[215] <=32'h38A218DF;
	Vec_Delta[216] <=32'h391AA60A;
	Vec_Delta[217] <=32'h39010C70;
	Vec_Delta[218] <=32'h38DD8696;
	Vec_Delta[219] <=32'h38C218DF;
	Vec_Delta[220] <=32'h39343FA3;
	Vec_Delta[221] <=32'h391661C5;
	Vec_Delta[222] <=32'h39010C70;
	Vec_Delta[223] <=32'h38E218DF;
	Vec_Delta[224] <=32'h3850FE8B;
	Vec_Delta[225] <=32'h382EDC69;
	Vec_Delta[226] <=32'h38167AE3;
	Vec_Delta[227] <=32'h380431BE;
	Vec_Delta[228] <=32'h388218DF;
	Vec_Delta[229] <=32'h38598714;
	Vec_Delta[230] <=32'h383B0D2C;
	Vec_Delta[231] <=32'h382431BE;
	Vec_Delta[232] <=32'h389BB279;
	Vec_Delta[233] <=32'h388218DF;
	Vec_Delta[234] <=32'h385F9F75;
	Vec_Delta[235] <=32'h384431BE;
	Vec_Delta[236] <=32'h38B54C13;
	Vec_Delta[237] <=32'h38976E35;
	Vec_Delta[238] <=32'h388218DF;
	Vec_Delta[239] <=32'h386431BE;
	Vec_Delta[240] <=32'h37D53049;
	Vec_Delta[241] <=32'h37B30E27;
	Vec_Delta[242] <=32'h379AACA1;
	Vec_Delta[243] <=32'h3788637C;
	Vec_Delta[244] <=32'h380431BE;
	Vec_Delta[245] <=32'h37DDB8D2;
	Vec_Delta[246] <=32'h37BF3EEA;
	Vec_Delta[247] <=32'h37A8637C;
	Vec_Delta[248] <=32'h381DCB58;
	Vec_Delta[249] <=32'h380431BE;
	Vec_Delta[250] <=32'h37E3D133;
	Vec_Delta[251] <=32'h37C8637C;
	Vec_Delta[252] <=32'h383764F2;
	Vec_Delta[253] <=32'h38198714;
	Vec_Delta[254] <=32'h380431BE;
	Vec_Delta[255] <=32'h37E8637C;
	
	//Theta circular vectoring
	Vec_Theta_Cir[0] <=32'h3F2CBBDD;
	Vec_Theta_Cir[1] <=32'h3F168762;
	Vec_Theta_Cir[2] <=32'h3F04E6CF;
	Vec_Theta_Cir[3] <=32'h3EED6353;
	Vec_Theta_Cir[4] <=32'h3F490FE3;
	Vec_Theta_Cir[5] <=32'h3F31DA68;
	Vec_Theta_Cir[6] <=32'h3F1EC8B7;
	Vec_Theta_Cir[7] <=32'h3F0F0069;
	Vec_Theta_Cir[8] <=32'h3F60455E;
	Vec_Theta_Cir[9] <=32'h3F490FE3;
	Vec_Theta_Cir[10] <=32'h3F356892;
	Vec_Theta_Cir[11] <=32'h3F24BC88;
	Vec_Theta_Cir[12] <=32'h3F735710;
	Vec_Theta_Cir[13] <=32'h3F5CB735;
	Vec_Theta_Cir[14] <=32'h3F490FE3;
	Vec_Theta_Cir[15] <=32'h3F380548;
	Vec_Theta_Cir[16] <=32'h3EC2D1D9;
	Vec_Theta_Cir[17] <=32'h3EA4BC9C;
	Vec_Theta_Cir[18] <=32'h3E8E7D6A;
	Vec_Theta_Cir[19] <=32'h3E7ADBEF;
	Vec_Theta_Cir[20] <=32'h3EED6354;
	Vec_Theta_Cir[21] <=32'h3ECA222D;
	Vec_Theta_Cir[22] <=32'h3EAFA0F3;
	Vec_Theta_Cir[23] <=32'h3E9B13D8;
	Vec_Theta_Cir[24] <=32'h3F0A58FB;
	Vec_Theta_Cir[25] <=32'h3EED6354;
	Vec_Theta_Cir[26] <=32'h3ECF4E17;
	Vec_Theta_Cir[27] <=32'h3EB7B0E8;
	Vec_Theta_Cir[28] <=32'h3F1C5895;
	Vec_Theta_Cir[29] <=32'h3F072FF0;
	Vec_Theta_Cir[30] <=32'h3EED6353;
	Vec_Theta_Cir[31] <=32'h3ED32793;
	Vec_Theta_Cir[32] <=32'h3E4A2251;
	Vec_Theta_Cir[33] <=32'h3E291CFE;
	Vec_Theta_Cir[34] <=32'h3E114DB8;
	Vec_Theta_Cir[35] <=32'h3DFEAE59;
	Vec_Theta_Cir[36] <=32'h3E7ADBF0;
	Vec_Theta_Cir[37] <=32'h3E52536C;
	Vec_Theta_Cir[38] <=32'h3E34F36C;
	Vec_Theta_Cir[39] <=32'h3E1EB7B9;
	Vec_Theta_Cir[40] <=32'h3E9539F2;
	Vec_Theta_Cir[41] <=32'h3E7ADBF0;
	Vec_Theta_Cir[42] <=32'h3E58291A;
	Vec_Theta_Cir[43] <=32'h3E3DCC1B;
	Vec_Theta_Cir[44] <=32'h3EAC60C3;
	Vec_Theta_Cir[45] <=32'h3E914D95;
	Vec_Theta_Cir[46] <=32'h3E7ADBF0;
	Vec_Theta_Cir[47] <=32'h3E5C86FB;
	Vec_Theta_Cir[48] <=32'h3DCC1F9A;
	Vec_Theta_Cir[49] <=32'h3DAA4679;
	Vec_Theta_Cir[50] <=32'h3D920A2C;
	Vec_Theta_Cir[51] <=32'h3D7FABEA;
	Vec_Theta_Cir[52] <=32'h3DFEAE5A;
	Vec_Theta_Cir[53] <=32'h3DD49199;
	Vec_Theta_Cir[54] <=32'h3DB66026;
	Vec_Theta_Cir[55] <=32'h3D9FAD7E;
	Vec_Theta_Cir[56] <=32'h3E1876DD;
	Vec_Theta_Cir[57] <=32'h3DFEAE5A;
	Vec_Theta_Cir[58] <=32'h3DDA98C1;
	Vec_Theta_Cir[59] <=32'h3DBF7146;
	Vec_Theta_Cir[60] <=32'h3E316792;
	Vec_Theta_Cir[61] <=32'h3E1449FC;
	Vec_Theta_Cir[62] <=32'h3DFEAE5A;
	Vec_Theta_Cir[63] <=32'h3DDF1D7B;
	Vec_Theta_Cir[64] <=32'h3D4CA239;
	Vec_Theta_Cir[65] <=32'h3D2A9275;
	Vec_Theta_Cir[66] <=32'h3D123A48;
	Vec_Theta_Cir[67] <=32'h3CFFECC7;
	Vec_Theta_Cir[68] <=32'h3D7FABEA;
	Vec_Theta_Cir[69] <=32'h3D552514;
	Vec_Theta_Cir[70] <=32'h3D36BD6A;
	Vec_Theta_Cir[71] <=32'h3D1FEC3C;
	Vec_Theta_Cir[72] <=32'h3D9950A5;
	Vec_Theta_Cir[73] <=32'h3D7FABEA;
	Vec_Theta_Cir[74] <=32'h3D5B391E;
	Vec_Theta_Cir[75] <=32'h3D3FDD18;
	Vec_Theta_Cir[76] <=32'h3DB2BF2E;
	Vec_Theta_Cir[77] <=32'h3D951251;
	Vec_Theta_Cir[78] <=32'h3D7FABEA;
	Vec_Theta_Cir[79] <=32'h3D5FC7FC;
	Vec_Theta_Cir[80] <=32'h3CCCC3FB;
	Vec_Theta_Cir[81] <=32'h3CAAA672;
	Vec_Theta_Cir[82] <=32'h3C924743;
	Vec_Theta_Cir[83] <=32'h3C7FFEDD;
	Vec_Theta_Cir[84] <=32'h3CFFECC7;
	Vec_Theta_Cir[85] <=32'h3CD54B17;
	Vec_Theta_Cir[86] <=32'h3CB6D5C1;
	Vec_Theta_Cir[87] <=32'h3C9FFCE4;
	Vec_Theta_Cir[88] <=32'h3D19883C;
	Vec_Theta_Cir[89] <=32'h3CFFECC7;
	Vec_Theta_Cir[90] <=32'h3CDB6262;
	Vec_Theta_Cir[91] <=32'h3CBFF91A;
	Vec_Theta_Cir[92] <=32'h3D331703;
	Vec_Theta_Cir[93] <=32'h3D154575;
	Vec_Theta_Cir[94] <=32'h3CFFECC7;
	Vec_Theta_Cir[95] <=32'h3CDFF3D0;
	Vec_Theta_Cir[96] <=32'h3C4CCE44;
	Vec_Theta_Cir[97] <=32'h3C2AAD48;
	Vec_Theta_Cir[98] <=32'h3C124C58;
	Vec_Theta_Cir[99] <=32'h3C000387;
	Vec_Theta_Cir[100] <=32'h3C7FFEDD;
	Vec_Theta_Cir[101] <=32'h3C555671;
	Vec_Theta_Cir[102] <=32'h3C36DDAE;
	Vec_Theta_Cir[103] <=32'h3C2002E4;
	Vec_Theta_Cir[104] <=32'h3C999717;
	Vec_Theta_Cir[105] <=32'h3C7FFEDD;
	Vec_Theta_Cir[106] <=32'h3C5B6E8D;
	Vec_Theta_Cir[107] <=32'h3C4001F2;
	Vec_Theta_Cir[108] <=32'h3CB32DFC;
	Vec_Theta_Cir[109] <=32'h3C955332;
	Vec_Theta_Cir[110] <=32'h3C7FFEDD;
	Vec_Theta_Cir[111] <=32'h3C60009F;
	Vec_Theta_Cir[112] <=32'h3BCCD482;
	Vec_Theta_Cir[113] <=32'h3BAAB2A9;
	Vec_Theta_Cir[114] <=32'h3B925148;
	Vec_Theta_Cir[115] <=32'h3B800839;
	Vec_Theta_Cir[116] <=32'h3C000387;
	Vec_Theta_Cir[117] <=32'h3BD55CF4;
	Vec_Theta_Cir[118] <=32'h3BB6E355;
	Vec_Theta_Cir[119] <=32'h3BA00810;
	Vec_Theta_Cir[120] <=32'h3C199CA5;
	Vec_Theta_Cir[121] <=32'h3C000387;
	Vec_Theta_Cir[122] <=32'h3BDB7544;
	Vec_Theta_Cir[123] <=32'h3BC007D4;
	Vec_Theta_Cir[124] <=32'h3C333591;
	Vec_Theta_Cir[125] <=32'h3C155878;
	Vec_Theta_Cir[126] <=32'h3C000387;
	Vec_Theta_Cir[127] <=32'h3BE0077F;
	Vec_Theta_Cir[128] <=32'h3B4CDD69;
	Vec_Theta_Cir[129] <=32'h3B2ABB59;
	Vec_Theta_Cir[130] <=32'h3B1259DC;
	Vec_Theta_Cir[131] <=32'h3B0010BC;
	Vec_Theta_Cir[132] <=32'h3B800839;
	Vec_Theta_Cir[133] <=32'h3B5565EB;
	Vec_Theta_Cir[134] <=32'h3B36EC16;
	Vec_Theta_Cir[135] <=32'h3B2010B2;
	Vec_Theta_Cir[136] <=32'h3B99A1B4;
	Vec_Theta_Cir[137] <=32'h3B800839;
	Vec_Theta_Cir[138] <=32'h3B5B7E49;
	Vec_Theta_Cir[139] <=32'h3B4010A3;
	Vec_Theta_Cir[140] <=32'h3BB33B22;
	Vec_Theta_Cir[141] <=32'h3B955D75;
	Vec_Theta_Cir[142] <=32'h3B800839;
	Vec_Theta_Cir[143] <=32'h3B60108E;
	Vec_Theta_Cir[144] <=32'h3ACCEE51;
	Vec_Theta_Cir[145] <=32'h3AAACC33;
	Vec_Theta_Cir[146] <=32'h3A926AAF;
	Vec_Theta_Cir[147] <=32'h3A80218B;
	Vec_Theta_Cir[148] <=32'h3B0010BD;
	Vec_Theta_Cir[149] <=32'h3AD576D8;
	Vec_Theta_Cir[150] <=32'h3AB6FCF4;
	Vec_Theta_Cir[151] <=32'h3AA02189;
	Vec_Theta_Cir[152] <=32'h3B19AA4F;
	Vec_Theta_Cir[153] <=32'h3B0010BC;
	Vec_Theta_Cir[154] <=32'h3ADB8F38;
	Vec_Theta_Cir[155] <=32'h3AC02185;
	Vec_Theta_Cir[156] <=32'h3B3343DD;
	Vec_Theta_Cir[157] <=32'h3B15660C;
	Vec_Theta_Cir[158] <=32'h3B0010BC;
	Vec_Theta_Cir[159] <=32'h3AE02180;
	Vec_Theta_Cir[160] <=32'h3A4D0FE7;
	Vec_Theta_Cir[161] <=32'h3A2AEDC5;
	Vec_Theta_Cir[162] <=32'h3A128C40;
	Vec_Theta_Cir[163] <=32'h3A00431B;
	Vec_Theta_Cir[164] <=32'h3A80218C;
	Vec_Theta_Cir[165] <=32'h3A55986F;
	Vec_Theta_Cir[166] <=32'h3A371E88;
	Vec_Theta_Cir[167] <=32'h3A20431B;
	Vec_Theta_Cir[168] <=32'h3A99BB23;
	Vec_Theta_Cir[169] <=32'h3A80218B;
	Vec_Theta_Cir[170] <=32'h3A5BB0D0;
	Vec_Theta_Cir[171] <=32'h3A40431A;
	Vec_Theta_Cir[172] <=32'h3AB354BA;
	Vec_Theta_Cir[173] <=32'h3A9576DF;
	Vec_Theta_Cir[174] <=32'h3A80218B;
	Vec_Theta_Cir[175] <=32'h3A604319;
	Vec_Theta_Cir[176] <=32'h39CD5305;
	Vec_Theta_Cir[177] <=32'h39AB30E2;
	Vec_Theta_Cir[178] <=32'h3992CF5C;
	Vec_Theta_Cir[179] <=32'h39808638;
	Vec_Theta_Cir[180] <=32'h3A00431B;
	Vec_Theta_Cir[181] <=32'h39D5DB8D;
	Vec_Theta_Cir[182] <=32'h39B761A5;
	Vec_Theta_Cir[183] <=32'h39A08638;
	Vec_Theta_Cir[184] <=32'h3A19DCB5;
	Vec_Theta_Cir[185] <=32'h3A00431B;
	Vec_Theta_Cir[186] <=32'h39DBF3EE;
	Vec_Theta_Cir[187] <=32'h39C08637;
	Vec_Theta_Cir[188] <=32'h3A33764E;
	Vec_Theta_Cir[189] <=32'h3A159870;
	Vec_Theta_Cir[190] <=32'h3A00431B;
	Vec_Theta_Cir[191] <=32'h39E08637;
	Vec_Theta_Cir[192] <=32'h394DD93D;
	Vec_Theta_Cir[193] <=32'h392BB71A;
	Vec_Theta_Cir[194] <=32'h39135594;
	Vec_Theta_Cir[195] <=32'h39010C6F;
	Vec_Theta_Cir[196] <=32'h39808638;
	Vec_Theta_Cir[197] <=32'h395661C5;
	Vec_Theta_Cir[198] <=32'h3937E7DD;
	Vec_Theta_Cir[199] <=32'h39210C70;
	Vec_Theta_Cir[200] <=32'h399A1FD2;
	Vec_Theta_Cir[201] <=32'h39808638;
	Vec_Theta_Cir[202] <=32'h395C7A27;
	Vec_Theta_Cir[203] <=32'h39410C70;
	Vec_Theta_Cir[204] <=32'h39B3B96B;
	Vec_Theta_Cir[205] <=32'h3995DB8D;
	Vec_Theta_Cir[206] <=32'h39808638;
	Vec_Theta_Cir[207] <=32'h39610C70;
	Vec_Theta_Cir[208] <=32'h38CEE5AC;
	Vec_Theta_Cir[209] <=32'h38ACC38A;
	Vec_Theta_Cir[210] <=32'h38946204;
	Vec_Theta_Cir[211] <=32'h388218DF;
	Vec_Theta_Cir[212] <=32'h39010C70;
	Vec_Theta_Cir[213] <=32'h38D76E35;
	Vec_Theta_Cir[214] <=32'h38B8F44D;
	Vec_Theta_Cir[215] <=32'h38A218DF;
	Vec_Theta_Cir[216] <=32'h391AA609;
	Vec_Theta_Cir[217] <=32'h39010C70;
	Vec_Theta_Cir[218] <=32'h38DD8696;
	Vec_Theta_Cir[219] <=32'h38C218DF;
	Vec_Theta_Cir[220] <=32'h39343FA3;
	Vec_Theta_Cir[221] <=32'h391661C5;
	Vec_Theta_Cir[222] <=32'h39010C70;
	Vec_Theta_Cir[223] <=32'h38E218DF;
	Vec_Theta_Cir[224] <=32'h3850FE8B;
	Vec_Theta_Cir[225] <=32'h382EDC69;
	Vec_Theta_Cir[226] <=32'h38167AE3;
	Vec_Theta_Cir[227] <=32'h380431BE;
	Vec_Theta_Cir[228] <=32'h388218DF;
	Vec_Theta_Cir[229] <=32'h38598714;
	Vec_Theta_Cir[230] <=32'h383B0D2C;
	Vec_Theta_Cir[231] <=32'h382431BE;
	Vec_Theta_Cir[232] <=32'h389BB279;
	Vec_Theta_Cir[233] <=32'h388218DF;
	Vec_Theta_Cir[234] <=32'h385F9F75;
	Vec_Theta_Cir[235] <=32'h384431BE;
	Vec_Theta_Cir[236] <=32'h38B54C13;
	Vec_Theta_Cir[237] <=32'h38976E35;
	Vec_Theta_Cir[238] <=32'h388218DF;
	Vec_Theta_Cir[239] <=32'h386431BE;
	Vec_Theta_Cir[240] <=32'h37D53049;
	Vec_Theta_Cir[241] <=32'h37B30E27;
	Vec_Theta_Cir[242] <=32'h379AACA1;
	Vec_Theta_Cir[243] <=32'h3788637C;
	Vec_Theta_Cir[244] <=32'h380431BE;
	Vec_Theta_Cir[245] <=32'h37DDB8D2;
	Vec_Theta_Cir[246] <=32'h37BF3EEA;
	Vec_Theta_Cir[247] <=32'h37A8637C;
	Vec_Theta_Cir[248] <=32'h381DCB58;
	Vec_Theta_Cir[249] <=32'h380431BE;
	Vec_Theta_Cir[250] <=32'h37E3D133;
	Vec_Theta_Cir[251] <=32'h37C8637C;
	Vec_Theta_Cir[252] <=32'h383764F2;
	Vec_Theta_Cir[253] <=32'h38198714;
	Vec_Theta_Cir[254] <=32'h380431BE;
	Vec_Theta_Cir[255] <=32'h37E8637C;
	
	//Theta vectoring hyperbolic
	Vec_Theta_Hyper[0] <=32'h3F8C9F6C;
	Vec_Theta_Hyper[1] <=32'h3F4E022F;
	Vec_Theta_Hyper[2] <=32'h3F264F01;
	Vec_Theta_Hyper[3] <=32'h3F0C9F6A;
	Vec_Theta_Hyper[4] <=32'h40E82375;
	Vec_Theta_Hyper[5] <=32'h3F99773B;
	Vec_Theta_Hyper[6] <=32'h3F655883;
	Vec_Theta_Hyper[7] <=32'h3F3BB10B;
	Vec_Theta_Hyper[8] <=32'h40E82375;
	Vec_Theta_Hyper[9] <=32'h40E82375;
	Vec_Theta_Hyper[10] <=32'h3FA42842;
	Vec_Theta_Hyper[11] <=32'h3F7913BD;
	Vec_Theta_Hyper[12] <=32'h40E82375;
	Vec_Theta_Hyper[13] <=32'h40E82375;
	Vec_Theta_Hyper[14] <=32'h40E82375;
	Vec_Theta_Hyper[15] <=32'h3FAD50D7;
	Vec_Theta_Hyper[16] <=32'h3ED8E8AC;
	Vec_Theta_Hyper[17] <=32'h3EB1723E;
	Vec_Theta_Hyper[18] <=32'h3E967955;
	Vec_Theta_Hyper[19] <=32'h3E82C59C;
	Vec_Theta_Hyper[20] <=32'h3F0C9F6B;
	Vec_Theta_Hyper[21] <=32'h3EE32677;
	Vec_Theta_Hyper[22] <=32'h3EBF4998;
	Vec_Theta_Hyper[23] <=32'h3EA58981;
	Vec_Theta_Hyper[24] <=32'h3F317233;
	Vec_Theta_Hyper[25] <=32'h3F0C9F6B;
	Vec_Theta_Hyper[26] <=32'h3EEA9231;
	Vec_Theta_Hyper[27] <=32'h3EC9D87F;
	Vec_Theta_Hyper[28] <=32'h3F5E078B;
	Vec_Theta_Hyper[29] <=32'h3F2AE16B;
	Vec_Theta_Hyper[30] <=32'h3F0C9F6A;
	Vec_Theta_Hyper[31] <=32'h3EF0329A;
	Vec_Theta_Hyper[32] <=32'h3E4F9966;
	Vec_Theta_Hyper[33] <=32'h3E2C465C;
	Vec_Theta_Hyper[34] <=32'h3E134B55;
	Vec_Theta_Hyper[35] <=32'h3E00AC8D;
	Vec_Theta_Hyper[36] <=32'h3E82C59C;
	Vec_Theta_Hyper[37] <=32'h3E5880F8;
	Vec_Theta_Hyper[38] <=32'h3E38D703;
	Vec_Theta_Hyper[39] <=32'h3E215292;
	Vec_Theta_Hyper[40] <=32'h3E9E7980;
	Vec_Theta_Hyper[41] <=32'h3E82C59C;
	Vec_Theta_Hyper[42] <=32'h3E5EE249;
	Vec_Theta_Hyper[43] <=32'h3E424CBD;
	Vec_Theta_Hyper[44] <=32'h3EBB1B99;
	Vec_Theta_Hyper[45] <=32'h3E99CC76;
	Vec_Theta_Hyper[46] <=32'h3E82C59C;
	Vec_Theta_Hyper[47] <=32'h3E63AE23;
	Vec_Theta_Hyper[48] <=32'h3DCD7D27;
	Vec_Theta_Hyper[49] <=32'h3DAB10C1;
	Vec_Theta_Hyper[50] <=32'h3D92898E;
	Vec_Theta_Hyper[51] <=32'h3D802B4B;
	Vec_Theta_Hyper[52] <=32'h3E00AC8D;
	Vec_Theta_Hyper[53] <=32'h3DD61CB1;
	Vec_Theta_Hyper[54] <=32'h3DB758F3;
	Vec_Theta_Hyper[55] <=32'h3DA0542B;
	Vec_Theta_Hyper[56] <=32'h3E1AC4D4;
	Vec_Theta_Hyper[57] <=32'h3E00AC8D;
	Vec_Theta_Hyper[58] <=32'h3DDC46B1;
	Vec_Theta_Hyper[59] <=32'h3DC0914B;
	Vec_Theta_Hyper[60] <=32'h3E351095;
	Vec_Theta_Hyper[61] <=32'h3E166820;
	Vec_Theta_Hyper[62] <=32'h3E00AC8D;
	Vec_Theta_Hyper[63] <=32'h3DE0E6DB;
	Vec_Theta_Hyper[64] <=32'h3D4CF99C;
	Vec_Theta_Hyper[65] <=32'h3D2AC507;
	Vec_Theta_Hyper[66] <=32'h3D125A21;
	Vec_Theta_Hyper[67] <=32'h3D000BB9;
	Vec_Theta_Hyper[68] <=32'h3D802B4B;
	Vec_Theta_Hyper[69] <=32'h3D5587DA;
	Vec_Theta_Hyper[70] <=32'h3D36FB9E;
	Vec_Theta_Hyper[71] <=32'h3D2015E7;
	Vec_Theta_Hyper[72] <=32'h3D99E41B;
	Vec_Theta_Hyper[73] <=32'h3D802B4B;
	Vec_Theta_Hyper[74] <=32'h3D5BA499;
	Vec_Theta_Hyper[75] <=32'h3D402519;
	Vec_Theta_Hyper[76] <=32'h3DB3A959;
	Vec_Theta_Hyper[77] <=32'h3D9599D5;
	Vec_Theta_Hyper[78] <=32'h3D802B4B;
	Vec_Theta_Hyper[79] <=32'h3D603A53;
	Vec_Theta_Hyper[80] <=32'h3CCCD9D4;
	Vec_Theta_Hyper[81] <=32'h3CAAB317;
	Vec_Theta_Hyper[82] <=32'h3C924F39;
	Vec_Theta_Hyper[83] <=32'h3C8004C4;
	Vec_Theta_Hyper[84] <=32'h3D000BB9;
	Vec_Theta_Hyper[85] <=32'h3CD563C9;
	Vec_Theta_Hyper[86] <=32'h3CB6E54E;
	Vec_Theta_Hyper[87] <=32'h3CA0074F;
	Vec_Theta_Hyper[88] <=32'h3D19AD19;
	Vec_Theta_Hyper[89] <=32'h3D000BB9;
	Vec_Theta_Hyper[90] <=32'h3CDB7D41;
	Vec_Theta_Hyper[91] <=32'h3CC00B1A;
	Vec_Theta_Hyper[92] <=32'h3D33518E;
	Vec_Theta_Hyper[93] <=32'h3D156756;
	Vec_Theta_Hyper[94] <=32'h3D000BB9;
	Vec_Theta_Hyper[95] <=32'h3CE01066;
	Vec_Theta_Hyper[96] <=32'h3C4CD3BB;
	Vec_Theta_Hyper[97] <=32'h3C2AB071;
	Vec_Theta_Hyper[98] <=32'h3C124E55;
	Vec_Theta_Hyper[99] <=32'h3C0004DC;
	Vec_Theta_Hyper[100] <=32'h3C8004C4;
	Vec_Theta_Hyper[101] <=32'h3C555C9E;
	Vec_Theta_Hyper[102] <=32'h3C36E192;
	Vec_Theta_Hyper[103] <=32'h3C20057F;
	Vec_Theta_Hyper[104] <=32'h3C99A04F;
	Vec_Theta_Hyper[105] <=32'h3C8004C4;
	Vec_Theta_Hyper[106] <=32'h3C5B7545;
	Vec_Theta_Hyper[107] <=32'h3C400672;
	Vec_Theta_Hyper[108] <=32'h3CB33C9F;
	Vec_Theta_Hyper[109] <=32'h3C955BAB;
	Vec_Theta_Hyper[110] <=32'h3C8004C4;
	Vec_Theta_Hyper[111] <=32'h3C6007C5;
	Vec_Theta_Hyper[112] <=32'h3BCCD5E0;
	Vec_Theta_Hyper[113] <=32'h3BAAB374;
	Vec_Theta_Hyper[114] <=32'h3B9251C8;
	Vec_Theta_Hyper[115] <=32'h3B80088E;
	Vec_Theta_Hyper[116] <=32'h3C0004DD;
	Vec_Theta_Hyper[117] <=32'h3BD55E7F;
	Vec_Theta_Hyper[118] <=32'h3BB6E44E;
	Vec_Theta_Hyper[119] <=32'h3BA008B7;
	Vec_Theta_Hyper[120] <=32'h3C199EF3;
	Vec_Theta_Hyper[121] <=32'h3C0004DD;
	Vec_Theta_Hyper[122] <=32'h3BDB76F2;
	Vec_Theta_Hyper[123] <=32'h3BC008F4;
	Vec_Theta_Hyper[124] <=32'h3C33393A;
	Vec_Theta_Hyper[125] <=32'h3C155A96;
	Vec_Theta_Hyper[126] <=32'h3C0004DD;
	Vec_Theta_Hyper[127] <=32'h3BE00949;
	Vec_Theta_Hyper[128] <=32'h3B4CDDC0;
	Vec_Theta_Hyper[129] <=32'h3B2ABB8B;
	Vec_Theta_Hyper[130] <=32'h3B1259FC;
	Vec_Theta_Hyper[131] <=32'h3B0010D2;
	Vec_Theta_Hyper[132] <=32'h3B80088E;
	Vec_Theta_Hyper[133] <=32'h3B55664E;
	Vec_Theta_Hyper[134] <=32'h3B36EC54;
	Vec_Theta_Hyper[135] <=32'h3B2010DC;
	Vec_Theta_Hyper[136] <=32'h3B99A247;
	Vec_Theta_Hyper[137] <=32'h3B80088E;
	Vec_Theta_Hyper[138] <=32'h3B5B7EB4;
	Vec_Theta_Hyper[139] <=32'h3B4010EB;
	Vec_Theta_Hyper[140] <=32'h3BB33C0C;
	Vec_Theta_Hyper[141] <=32'h3B955DFD;
	Vec_Theta_Hyper[142] <=32'h3B80088E;
	Vec_Theta_Hyper[143] <=32'h3B601101;
	Vec_Theta_Hyper[144] <=32'h3ACCEE66;
	Vec_Theta_Hyper[145] <=32'h3AAACC3F;
	Vec_Theta_Hyper[146] <=32'h3A926AB7;
	Vec_Theta_Hyper[147] <=32'h3A802191;
	Vec_Theta_Hyper[148] <=32'h3B0010D2;
	Vec_Theta_Hyper[149] <=32'h3AD576F0;
	Vec_Theta_Hyper[150] <=32'h3AB6FD04;
	Vec_Theta_Hyper[151] <=32'h3AA02193;
	Vec_Theta_Hyper[152] <=32'h3B19AA73;
	Vec_Theta_Hyper[153] <=32'h3B0010D2;
	Vec_Theta_Hyper[154] <=32'h3ADB8F53;
	Vec_Theta_Hyper[155] <=32'h3AC02197;
	Vec_Theta_Hyper[156] <=32'h3B334418;
	Vec_Theta_Hyper[157] <=32'h3B15662E;
	Vec_Theta_Hyper[158] <=32'h3B0010D2;
	Vec_Theta_Hyper[159] <=32'h3AE0219D;
	Vec_Theta_Hyper[160] <=32'h3A4D0FEC;
	Vec_Theta_Hyper[161] <=32'h3A2AEDC9;
	Vec_Theta_Hyper[162] <=32'h3A128C42;
	Vec_Theta_Hyper[163] <=32'h3A00431D;
	Vec_Theta_Hyper[164] <=32'h3A802191;
	Vec_Theta_Hyper[165] <=32'h3A559875;
	Vec_Theta_Hyper[166] <=32'h3A371E8C;
	Vec_Theta_Hyper[167] <=32'h3A20431D;
	Vec_Theta_Hyper[168] <=32'h3A99BB2D;
	Vec_Theta_Hyper[169] <=32'h3A802191;
	Vec_Theta_Hyper[170] <=32'h3A5BB0D7;
	Vec_Theta_Hyper[171] <=32'h3A40431E;
	Vec_Theta_Hyper[172] <=32'h3AB354C9;
	Vec_Theta_Hyper[173] <=32'h3A9576E8;
	Vec_Theta_Hyper[174] <=32'h3A802191;
	Vec_Theta_Hyper[175] <=32'h3A604320;
	Vec_Theta_Hyper[176] <=32'h39CD5306;
	Vec_Theta_Hyper[177] <=32'h39AB30E3;
	Vec_Theta_Hyper[178] <=32'h3992CF5D;
	Vec_Theta_Hyper[179] <=32'h39808638;
	Vec_Theta_Hyper[180] <=32'h3A00431D;
	Vec_Theta_Hyper[181] <=32'h39D5DB8E;
	Vec_Theta_Hyper[182] <=32'h39B761A6;
	Vec_Theta_Hyper[183] <=32'h39A08638;
	Vec_Theta_Hyper[184] <=32'h3A19DCB7;
	Vec_Theta_Hyper[185] <=32'h3A00431D;
	Vec_Theta_Hyper[186] <=32'h39DBF3F0;
	Vec_Theta_Hyper[187] <=32'h39C08639;
	Vec_Theta_Hyper[188] <=32'h3A337652;
	Vec_Theta_Hyper[189] <=32'h3A159873;
	Vec_Theta_Hyper[190] <=32'h3A00431D;
	Vec_Theta_Hyper[191] <=32'h39E08639;
	Vec_Theta_Hyper[192] <=32'h394DD93D;
	Vec_Theta_Hyper[193] <=32'h392BB71B;
	Vec_Theta_Hyper[194] <=32'h39135594;
	Vec_Theta_Hyper[195] <=32'h39010C70;
	Vec_Theta_Hyper[196] <=32'h39808638;
	Vec_Theta_Hyper[197] <=32'h395661C6;
	Vec_Theta_Hyper[198] <=32'h3937E7DE;
	Vec_Theta_Hyper[199] <=32'h39210C70;
	Vec_Theta_Hyper[200] <=32'h399A1FD2;
	Vec_Theta_Hyper[201] <=32'h39808638;
	Vec_Theta_Hyper[202] <=32'h395C7A27;
	Vec_Theta_Hyper[203] <=32'h39410C70;
	Vec_Theta_Hyper[204] <=32'h39B3B96C;
	Vec_Theta_Hyper[205] <=32'h3995DB8E;
	Vec_Theta_Hyper[206] <=32'h39808638;
	Vec_Theta_Hyper[207] <=32'h39610C70;
	Vec_Theta_Hyper[208] <=32'h38CEE5AD;
	Vec_Theta_Hyper[209] <=32'h38ACC38A;
	Vec_Theta_Hyper[210] <=32'h38946204;
	Vec_Theta_Hyper[211] <=32'h388218DF;
	Vec_Theta_Hyper[212] <=32'h39010C70;
	Vec_Theta_Hyper[213] <=32'h38D76E35;
	Vec_Theta_Hyper[214] <=32'h38B8F44D;
	Vec_Theta_Hyper[215] <=32'h38A218DF;
	Vec_Theta_Hyper[216] <=32'h391AA60A;
	Vec_Theta_Hyper[217] <=32'h39010C70;
	Vec_Theta_Hyper[218] <=32'h38DD8696;
	Vec_Theta_Hyper[219] <=32'h38C218DF;
	Vec_Theta_Hyper[220] <=32'h39343FA3;
	Vec_Theta_Hyper[221] <=32'h391661C5;
	Vec_Theta_Hyper[222] <=32'h39010C70;
	Vec_Theta_Hyper[223] <=32'h38E218DF;
	Vec_Theta_Hyper[224] <=32'h3850FE8B;
	Vec_Theta_Hyper[225] <=32'h382EDC69;
	Vec_Theta_Hyper[226] <=32'h38167AE3;
	Vec_Theta_Hyper[227] <=32'h380431BE;
	Vec_Theta_Hyper[228] <=32'h388218DF;
	Vec_Theta_Hyper[229] <=32'h38598714;
	Vec_Theta_Hyper[230] <=32'h383B0D2C;
	Vec_Theta_Hyper[231] <=32'h382431BE;
	Vec_Theta_Hyper[232] <=32'h389BB279;
	Vec_Theta_Hyper[233] <=32'h388218DF;
	Vec_Theta_Hyper[234] <=32'h385F9F75;
	Vec_Theta_Hyper[235] <=32'h384431BE;
	Vec_Theta_Hyper[236] <=32'h38B54C13;
	Vec_Theta_Hyper[237] <=32'h38976E35;
	Vec_Theta_Hyper[238] <=32'h388218DF;
	Vec_Theta_Hyper[239] <=32'h386431BE;
	Vec_Theta_Hyper[240] <=32'h37D53049;
	Vec_Theta_Hyper[241] <=32'h37B30E27;
	Vec_Theta_Hyper[242] <=32'h379AACA1;
	Vec_Theta_Hyper[243] <=32'h3788637C;
	Vec_Theta_Hyper[244] <=32'h380431BE;
	Vec_Theta_Hyper[245] <=32'h37DDB8D2;
	Vec_Theta_Hyper[246] <=32'h37BF3EEA;
	Vec_Theta_Hyper[247] <=32'h37A8637C;
	Vec_Theta_Hyper[248] <=32'h381DCB58;
	Vec_Theta_Hyper[249] <=32'h380431BE;
	Vec_Theta_Hyper[250] <=32'h37E3D133;
	Vec_Theta_Hyper[251] <=32'h37C8637C;
	Vec_Theta_Hyper[252] <=32'h383764F2;
	Vec_Theta_Hyper[253] <=32'h38198714;
	Vec_Theta_Hyper[254] <=32'h380431BE;
	Vec_Theta_Hyper[255] <=32'h37E8637C;
	
	//Kappa vectoring hyperbolic
	Vec_Kappa_Hyper[0] <=32'h3FD5557A;
	Vec_Kappa_Hyper[1] <=32'h3FABBAF5;
	Vec_Kappa_Hyper[2] <=32'h3F9BF949;
	Vec_Kappa_Hyper[3] <=32'h3F93CD45;
	Vec_Kappa_Hyper[4] <=32'h4430C6D8;
	Vec_Kappa_Hyper[5] <=32'h3FE78FBB;
	Vec_Kappa_Hyper[6] <=32'h3FB6E544;
	Vec_Kappa_Hyper[7] <=32'h3FA3F8B2;
	Vec_Kappa_Hyper[8] <=32'h4430C6D8;
	Vec_Kappa_Hyper[9] <=32'h4430C6D8;
	Vec_Kappa_Hyper[10] <=32'h3FF881B0;
	Vec_Kappa_Hyper[11] <=32'h3FC184AA;
	Vec_Kappa_Hyper[12] <=32'h4430C6D8;
	Vec_Kappa_Hyper[13] <=32'h4430C6D8;
	Vec_Kappa_Hyper[14] <=32'h4430C6D8;
	Vec_Kappa_Hyper[15] <=32'h400432C9;
	Vec_Kappa_Hyper[16] <=32'h3F8BA8DA;
	Vec_Kappa_Hyper[17] <=32'h3F87C3BE;
	Vec_Kappa_Hyper[18] <=32'h3F859161;
	Vec_Kappa_Hyper[19] <=32'h3F8432AB;
	Vec_Kappa_Hyper[20] <=32'h3F93CD45;
	Vec_Kappa_Hyper[21] <=32'h3F8CCE16;
	Vec_Kappa_Hyper[22] <=32'h3F8909AC;
	Vec_Kappa_Hyper[23] <=32'h3F86BFA5;
	Vec_Kappa_Hyper[24] <=32'h3FA0000E;
	Vec_Kappa_Hyper[25] <=32'h3F93CD45;
	Vec_Kappa_Hyper[26] <=32'h3F8DAB90;
	Vec_Kappa_Hyper[27] <=32'h3F8A1385;
	Vec_Kappa_Hyper[28] <=32'h3FB33C76;
	Vec_Kappa_Hyper[29] <=32'h3F9D972A;
	Vec_Kappa_Hyper[30] <=32'h3F93CD45;
	Vec_Kappa_Hyper[31] <=32'h3F8E5892;
	Vec_Kappa_Hyper[32] <=32'h3F82A3B9;
	Vec_Kappa_Hyper[33] <=32'h3F81D0D6;
	Vec_Kappa_Hyper[34] <=32'h3F815398;
	Vec_Kappa_Hyper[35] <=32'h3F81030F;
	Vec_Kappa_Hyper[36] <=32'h3F8432AB;
	Vec_Kappa_Hyper[37] <=32'h3F82DF27;
	Vec_Kappa_Hyper[38] <=32'h3F82174E;
	Vec_Kappa_Hyper[39] <=32'h3F81977F;
	Vec_Kappa_Hyper[40] <=32'h3F862E39;
	Vec_Kappa_Hyper[41] <=32'h3F8432AB;
	Vec_Kappa_Hyper[42] <=32'h3F830B4A;
	Vec_Kappa_Hyper[43] <=32'h3F824FAB;
	Vec_Kappa_Hyper[44] <=32'h3F88A48F;
	Vec_Kappa_Hyper[45] <=32'h3F85D18B;
	Vec_Kappa_Hyper[46] <=32'h3F8432AB;
	Vec_Kappa_Hyper[47] <=32'h3F832D54;
	Vec_Kappa_Hyper[48] <=32'h3F80A519;
	Vec_Kappa_Hyper[49] <=32'h3F807264;
	Vec_Kappa_Hyper[50] <=32'h3F8053EE;
	Vec_Kappa_Hyper[51] <=32'h3F804034;
	Vec_Kappa_Hyper[52] <=32'h3F81030F;
	Vec_Kappa_Hyper[53] <=32'h3F80B341;
	Vec_Kappa_Hyper[54] <=32'h3F80836A;
	Vec_Kappa_Hyper[55] <=32'h3F80647A;
	Vec_Kappa_Hyper[56] <=32'h3F817700;
	Vec_Kappa_Hyper[57] <=32'h3F81030F;
	Vec_Kappa_Hyper[58] <=32'h3F80BDBC;
	Vec_Kappa_Hyper[59] <=32'h3F8090F9;
	Vec_Kappa_Hyper[60] <=32'h3F82019C;
	Vec_Kappa_Hyper[61] <=32'h3F81621F;
	Vec_Kappa_Hyper[62] <=32'h3F81030F;
	Vec_Kappa_Hyper[63] <=32'h3F80C5CB;
	Vec_Kappa_Hyper[64] <=32'h3F80290E;
	Vec_Kappa_Hyper[65] <=32'h3F801C7F;
	Vec_Kappa_Hyper[66] <=32'h3F8014EF;
	Vec_Kappa_Hyper[67] <=32'h3F801007;
	Vec_Kappa_Hyper[68] <=32'h3F804034;
	Vec_Kappa_Hyper[69] <=32'h3F802C8D;
	Vec_Kappa_Hyper[70] <=32'h3F8020B8;
	Vec_Kappa_Hyper[71] <=32'h3F80190B;
	Vec_Kappa_Hyper[72] <=32'h3F805C91;
	Vec_Kappa_Hyper[73] <=32'h3F804034;
	Vec_Kappa_Hyper[74] <=32'h3F802F23;
	Vec_Kappa_Hyper[75] <=32'h3F802413;
	Vec_Kappa_Hyper[76] <=32'h3F807E2F;
	Vec_Kappa_Hyper[77] <=32'h3F80577A;
	Vec_Kappa_Hyper[78] <=32'h3F804034;
	Vec_Kappa_Hyper[79] <=32'h3F803120;
	Vec_Kappa_Hyper[80] <=32'h3F800A43;
	Vec_Kappa_Hyper[81] <=32'h3F800721;
	Vec_Kappa_Hyper[82] <=32'h3F80053E;
	Vec_Kappa_Hyper[83] <=32'h3F800404;
	Vec_Kappa_Hyper[84] <=32'h3F801007;
	Vec_Kappa_Hyper[85] <=32'h3F800B22;
	Vec_Kappa_Hyper[86] <=32'h3F80082E;
	Vec_Kappa_Hyper[87] <=32'h3F800644;
	Vec_Kappa_Hyper[88] <=32'h3F801714;
	Vec_Kappa_Hyper[89] <=32'h3F801007;
	Vec_Kappa_Hyper[90] <=32'h3F800BC7;
	Vec_Kappa_Hyper[91] <=32'h3F800905;
	Vec_Kappa_Hyper[92] <=32'h3F801F6C;
	Vec_Kappa_Hyper[93] <=32'h3F8015D1;
	Vec_Kappa_Hyper[94] <=32'h3F801007;
	Vec_Kappa_Hyper[95] <=32'h3F800C46;
	Vec_Kappa_Hyper[96] <=32'h3F800293;
	Vec_Kappa_Hyper[97] <=32'h3F8001CB;
	Vec_Kappa_Hyper[98] <=32'h3F800152;
	Vec_Kappa_Hyper[99] <=32'h3F800104;
	Vec_Kappa_Hyper[100] <=32'h3F800404;
	Vec_Kappa_Hyper[101] <=32'h3F8002CB;
	Vec_Kappa_Hyper[102] <=32'h3F80020E;
	Vec_Kappa_Hyper[103] <=32'h3F800194;
	Vec_Kappa_Hyper[104] <=32'h3F8005C7;
	Vec_Kappa_Hyper[105] <=32'h3F800404;
	Vec_Kappa_Hyper[106] <=32'h3F8002F4;
	Vec_Kappa_Hyper[107] <=32'h3F800244;
	Vec_Kappa_Hyper[108] <=32'h3F8007DC;
	Vec_Kappa_Hyper[109] <=32'h3F800576;
	Vec_Kappa_Hyper[110] <=32'h3F800404;
	Vec_Kappa_Hyper[111] <=32'h3F800314;
	Vec_Kappa_Hyper[112] <=32'h3F8000A8;
	Vec_Kappa_Hyper[113] <=32'h3F800076;
	Vec_Kappa_Hyper[114] <=32'h3F800057;
	Vec_Kappa_Hyper[115] <=32'h3F800044;
	Vec_Kappa_Hyper[116] <=32'h3F800104;
	Vec_Kappa_Hyper[117] <=32'h3F8000B6;
	Vec_Kappa_Hyper[118] <=32'h3F800086;
	Vec_Kappa_Hyper[119] <=32'h3F800068;
	Vec_Kappa_Hyper[120] <=32'h3F800174;
	Vec_Kappa_Hyper[121] <=32'h3F800104;
	Vec_Kappa_Hyper[122] <=32'h3F8000C0;
	Vec_Kappa_Hyper[123] <=32'h3F800094;
	Vec_Kappa_Hyper[124] <=32'h3F8001FA;
	Vec_Kappa_Hyper[125] <=32'h3F800160;
	Vec_Kappa_Hyper[126] <=32'h3F800104;
	Vec_Kappa_Hyper[127] <=32'h3F8000C8;
	Vec_Kappa_Hyper[128] <=32'h3F80002D;
	Vec_Kappa_Hyper[129] <=32'h3F800020;
	Vec_Kappa_Hyper[130] <=32'h3F800019;
	Vec_Kappa_Hyper[131] <=32'h3F800014;
	Vec_Kappa_Hyper[132] <=32'h3F800044;
	Vec_Kappa_Hyper[133] <=32'h3F800030;
	Vec_Kappa_Hyper[134] <=32'h3F800024;
	Vec_Kappa_Hyper[135] <=32'h3F80001D;
	Vec_Kappa_Hyper[136] <=32'h3F800060;
	Vec_Kappa_Hyper[137] <=32'h3F800044;
	Vec_Kappa_Hyper[138] <=32'h3F800033;
	Vec_Kappa_Hyper[139] <=32'h3F800028;
	Vec_Kappa_Hyper[140] <=32'h3F800081;
	Vec_Kappa_Hyper[141] <=32'h3F80005B;
	Vec_Kappa_Hyper[142] <=32'h3F800044;
	Vec_Kappa_Hyper[143] <=32'h3F800035;
	Vec_Kappa_Hyper[144] <=32'h3F80000E;
	Vec_Kappa_Hyper[145] <=32'h3F80000B;
	Vec_Kappa_Hyper[146] <=32'h3F800009;
	Vec_Kappa_Hyper[147] <=32'h3F800008;
	Vec_Kappa_Hyper[148] <=32'h3F800014;
	Vec_Kappa_Hyper[149] <=32'h3F80000F;
	Vec_Kappa_Hyper[150] <=32'h3F80000C;
	Vec_Kappa_Hyper[151] <=32'h3F80000A;
	Vec_Kappa_Hyper[152] <=32'h3F80001B;
	Vec_Kappa_Hyper[153] <=32'h3F800014;
	Vec_Kappa_Hyper[154] <=32'h3F80000F;
	Vec_Kappa_Hyper[155] <=32'h3F80000D;
	Vec_Kappa_Hyper[156] <=32'h3F800023;
	Vec_Kappa_Hyper[157] <=32'h3F800019;
	Vec_Kappa_Hyper[158] <=32'h3F800014;
	Vec_Kappa_Hyper[159] <=32'h3F800010;
	Vec_Kappa_Hyper[160] <=32'h3F800006;
	Vec_Kappa_Hyper[161] <=32'h3F800005;
	Vec_Kappa_Hyper[162] <=32'h3F800005;
	Vec_Kappa_Hyper[163] <=32'h3F800005;
	Vec_Kappa_Hyper[164] <=32'h3F800008;
	Vec_Kappa_Hyper[165] <=32'h3F800006;
	Vec_Kappa_Hyper[166] <=32'h3F800006;
	Vec_Kappa_Hyper[167] <=32'h3F800005;
	Vec_Kappa_Hyper[168] <=32'h3F800009;
	Vec_Kappa_Hyper[169] <=32'h3F800008;
	Vec_Kappa_Hyper[170] <=32'h3F800007;
	Vec_Kappa_Hyper[171] <=32'h3F800006;
	Vec_Kappa_Hyper[172] <=32'h3F80000C;
	Vec_Kappa_Hyper[173] <=32'h3F800009;
	Vec_Kappa_Hyper[174] <=32'h3F800008;
	Vec_Kappa_Hyper[175] <=32'h3F800007;
	Vec_Kappa_Hyper[176] <=32'h3F800004;
	Vec_Kappa_Hyper[177] <=32'h3F800004;
	Vec_Kappa_Hyper[178] <=32'h3F800004;
	Vec_Kappa_Hyper[179] <=32'h3F800004;
	Vec_Kappa_Hyper[180] <=32'h3F800005;
	Vec_Kappa_Hyper[181] <=32'h3F800004;
	Vec_Kappa_Hyper[182] <=32'h3F800004;
	Vec_Kappa_Hyper[183] <=32'h3F800004;
	Vec_Kappa_Hyper[184] <=32'h3F800005;
	Vec_Kappa_Hyper[185] <=32'h3F800005;
	Vec_Kappa_Hyper[186] <=32'h3F800004;
	Vec_Kappa_Hyper[187] <=32'h3F800004;
	Vec_Kappa_Hyper[188] <=32'h3F800006;
	Vec_Kappa_Hyper[189] <=32'h3F800005;
	Vec_Kappa_Hyper[190] <=32'h3F800005;
	Vec_Kappa_Hyper[191] <=32'h3F800004;
	Vec_Kappa_Hyper[192] <=32'h3F800004;
	Vec_Kappa_Hyper[193] <=32'h3F800004;
	Vec_Kappa_Hyper[194] <=32'h3F800004;
	Vec_Kappa_Hyper[195] <=32'h3F800004;
	Vec_Kappa_Hyper[196] <=32'h3F800004;
	Vec_Kappa_Hyper[197] <=32'h3F800004;
	Vec_Kappa_Hyper[198] <=32'h3F800004;
	Vec_Kappa_Hyper[199] <=32'h3F800004;
	Vec_Kappa_Hyper[200] <=32'h3F800004;
	Vec_Kappa_Hyper[201] <=32'h3F800004;
	Vec_Kappa_Hyper[202] <=32'h3F800004;
	Vec_Kappa_Hyper[203] <=32'h3F800004;
	Vec_Kappa_Hyper[204] <=32'h3F800004;
	Vec_Kappa_Hyper[205] <=32'h3F800004;
	Vec_Kappa_Hyper[206] <=32'h3F800004;
	Vec_Kappa_Hyper[207] <=32'h3F800004;
	Vec_Kappa_Hyper[208] <=32'h3F800004;
	Vec_Kappa_Hyper[209] <=32'h3F800004;
	Vec_Kappa_Hyper[210] <=32'h3F800004;
	Vec_Kappa_Hyper[211] <=32'h3F800004;
	Vec_Kappa_Hyper[212] <=32'h3F800004;
	Vec_Kappa_Hyper[213] <=32'h3F800004;
	Vec_Kappa_Hyper[214] <=32'h3F800004;
	Vec_Kappa_Hyper[215] <=32'h3F800004;
	Vec_Kappa_Hyper[216] <=32'h3F800004;
	Vec_Kappa_Hyper[217] <=32'h3F800004;
	Vec_Kappa_Hyper[218] <=32'h3F800004;
	Vec_Kappa_Hyper[219] <=32'h3F800004;
	Vec_Kappa_Hyper[220] <=32'h3F800004;
	Vec_Kappa_Hyper[221] <=32'h3F800004;
	Vec_Kappa_Hyper[222] <=32'h3F800004;
	Vec_Kappa_Hyper[223] <=32'h3F800004;
	Vec_Kappa_Hyper[224] <=32'h3F800004;
	Vec_Kappa_Hyper[225] <=32'h3F800004;
	Vec_Kappa_Hyper[226] <=32'h3F800004;
	Vec_Kappa_Hyper[227] <=32'h3F800004;
	Vec_Kappa_Hyper[228] <=32'h3F800004;
	Vec_Kappa_Hyper[229] <=32'h3F800004;
	Vec_Kappa_Hyper[230] <=32'h3F800004;
	Vec_Kappa_Hyper[231] <=32'h3F800004;
	Vec_Kappa_Hyper[232] <=32'h3F800004;
	Vec_Kappa_Hyper[233] <=32'h3F800004;
	Vec_Kappa_Hyper[234] <=32'h3F800004;
	Vec_Kappa_Hyper[235] <=32'h3F800004;
	Vec_Kappa_Hyper[236] <=32'h3F800004;
	Vec_Kappa_Hyper[237] <=32'h3F800004;
	Vec_Kappa_Hyper[238] <=32'h3F800004;
	Vec_Kappa_Hyper[239] <=32'h3F800004;
	Vec_Kappa_Hyper[240] <=32'h3F800004;
	Vec_Kappa_Hyper[241] <=32'h3F800004;
	Vec_Kappa_Hyper[242] <=32'h3F800004;
	Vec_Kappa_Hyper[243] <=32'h3F800004;
	Vec_Kappa_Hyper[244] <=32'h3F800004;
	Vec_Kappa_Hyper[245] <=32'h3F800004;
	Vec_Kappa_Hyper[246] <=32'h3F800004;
	Vec_Kappa_Hyper[247] <=32'h3F800004;
	Vec_Kappa_Hyper[248] <=32'h3F800004;
	Vec_Kappa_Hyper[249] <=32'h3F800004;
	Vec_Kappa_Hyper[250] <=32'h3F800004;
	Vec_Kappa_Hyper[251] <=32'h3F800004;
	Vec_Kappa_Hyper[252] <=32'h3F800004;
	Vec_Kappa_Hyper[253] <=32'h3F800004;
	Vec_Kappa_Hyper[254] <=32'h3F800004;
	Vec_Kappa_Hyper[255] <=32'h3F800004;
	
	//Kappa vectoring circular
	Vec_Kappa_Cir[0] <=32'h3F47E706;
	Vec_Kappa_Cir[1] <=32'h3F550141;
	Vec_Kappa_Cir[2] <=32'h3F5E4530;
	Vec_Kappa_Cir[3] <=32'h3F64F930;
	Vec_Kappa_Cir[4] <=32'h3F3504F5;
	Vec_Kappa_Cir[5] <=32'h3F44AA27;
	Vec_Kappa_Cir[6] <=32'h3F5050D7;
	Vec_Kappa_Cir[7] <=32'h3F59166C;
	Vec_Kappa_Cir[8] <=32'h3F23E322;
	Vec_Kappa_Cir[9] <=32'h3F3504F5;
	Vec_Kappa_Cir[10] <=32'h3F425EA5;
	Vec_Kappa_Cir[11] <=32'h3F4CCCCE;
	Vec_Kappa_Cir[12] <=32'h3F14CC09;
	Vec_Kappa_Cir[13] <=32'h3F269A45;
	Vec_Kappa_Cir[14] <=32'h3F3504F5;
	Vec_Kappa_Cir[15] <=32'h3F40A8DF;
	Vec_Kappa_Cir[16] <=32'h3F6DB0A8;
	Vec_Kappa_Cir[17] <=32'h3F72DCEC;
	Vec_Kappa_Cir[18] <=32'h3F762673;
	Vec_Kappa_Cir[19] <=32'h3F785B46;
	Vec_Kappa_Cir[20] <=32'h3F64F930;
	Vec_Kappa_Cir[21] <=32'h3F6C4EC7;
	Vec_Kappa_Cir[22] <=32'h3F711602;
	Vec_Kappa_Cir[23] <=32'h3F7458D0;
	Vec_Kappa_Cir[24] <=32'h3F5B84A9;
	Vec_Kappa_Cir[25] <=32'h3F64F930;
	Vec_Kappa_Cir[26] <=32'h3F6B4D19;
	Vec_Kappa_Cir[27] <=32'h3F6FB347;
	Vec_Kappa_Cir[28] <=32'h3F51B930;
	Vec_Kappa_Cir[29] <=32'h3F5D209E;
	Vec_Kappa_Cir[30] <=32'h3F64F930;
	Vec_Kappa_Cir[31] <=32'h3F6A894C;
	Vec_Kappa_Cir[32] <=32'h3F7B075A;
	Vec_Kappa_Cir[33] <=32'h3F7C8455;
	Vec_Kappa_Cir[34] <=32'h3F7D6D5A;
	Vec_Kappa_Cir[35] <=32'h3F7E05F2;
	Vec_Kappa_Cir[36] <=32'h3F785B46;
	Vec_Kappa_Cir[37] <=32'h3F7A9E7B;
	Vec_Kappa_Cir[38] <=32'h3F7C0377;
	Vec_Kappa_Cir[39] <=32'h3F7CEE61;
	Vec_Kappa_Cir[40] <=32'h3F75341E;
	Vec_Kappa_Cir[41] <=32'h3F785B46;
	Vec_Kappa_Cir[42] <=32'h3F7A5147;
	Vec_Kappa_Cir[43] <=32'h3F7B9D88;
	Vec_Kappa_Cir[44] <=32'h3F71A0B6;
	Vec_Kappa_Cir[45] <=32'h3F75C293;
	Vec_Kappa_Cir[46] <=32'h3F785B46;
	Vec_Kappa_Cir[47] <=32'h3F7A1623;
	Vec_Kappa_Cir[48] <=32'h3F7EBAC8;
	Vec_Kappa_Cir[49] <=32'h3F7F1DA6;
	Vec_Kappa_Cir[50] <=32'h3F7F597B;
	Vec_Kappa_Cir[51] <=32'h3F7F8067;
	Vec_Kappa_Cir[52] <=32'h3F7E05F2;
	Vec_Kappa_Cir[53] <=32'h3F7E9F56;
	Vec_Kappa_Cir[54] <=32'h3F7EFC5A;
	Vec_Kappa_Cir[55] <=32'h3F7F38F0;
	Vec_Kappa_Cir[56] <=32'h3F7D2AF4;
	Vec_Kappa_Cir[57] <=32'h3F7E05F2;
	Vec_Kappa_Cir[58] <=32'h3F7E8B12;
	Vec_Kappa_Cir[59] <=32'h3F7EE1E9;
	Vec_Kappa_Cir[60] <=32'h3F7C2AFA;
	Vec_Kappa_Cir[61] <=32'h3F7D520E;
	Vec_Kappa_Cir[62] <=32'h3F7E05F2;
	Vec_Kappa_Cir[63] <=32'h3F7E7B82;
	Vec_Kappa_Cir[64] <=32'h3F7FAE43;
	Vec_Kappa_Cir[65] <=32'h3F7FC737;
	Vec_Kappa_Cir[66] <=32'h3F7FD646;
	Vec_Kappa_Cir[67] <=32'h3F7FE00D;
	Vec_Kappa_Cir[68] <=32'h3F7F8067;
	Vec_Kappa_Cir[69] <=32'h3F7FA752;
	Vec_Kappa_Cir[70] <=32'h3F7FBED2;
	Vec_Kappa_Cir[71] <=32'h3F7FCE16;
	Vec_Kappa_Cir[72] <=32'h3F7F487B;
	Vec_Kappa_Cir[73] <=32'h3F7F8067;
	Vec_Kappa_Cir[74] <=32'h3F7FA230;
	Vec_Kappa_Cir[75] <=32'h3F7FB825;
	Vec_Kappa_Cir[76] <=32'h3F7F0694;
	Vec_Kappa_Cir[77] <=32'h3F7F527F;
	Vec_Kappa_Cir[78] <=32'h3F7F8067;
	Vec_Kappa_Cir[79] <=32'h3F7F9E3F;
	Vec_Kappa_Cir[80] <=32'h3F7FEB8F;
	Vec_Kappa_Cir[81] <=32'h3F7FF1D0;
	Vec_Kappa_Cir[82] <=32'h3F7FF595;
	Vec_Kappa_Cir[83] <=32'h3F7FF808;
	Vec_Kappa_Cir[84] <=32'h3F7FE00D;
	Vec_Kappa_Cir[85] <=32'h3F7FE9D1;
	Vec_Kappa_Cir[86] <=32'h3F7FEFB5;
	Vec_Kappa_Cir[87] <=32'h3F7FF388;
	Vec_Kappa_Cir[88] <=32'h3F7FD1FF;
	Vec_Kappa_Cir[89] <=32'h3F7FE00D;
	Vec_Kappa_Cir[90] <=32'h3F7FE888;
	Vec_Kappa_Cir[91] <=32'h3F7FEE09;
	Vec_Kappa_Cir[92] <=32'h3F7FC166;
	Vec_Kappa_Cir[93] <=32'h3F7FD484;
	Vec_Kappa_Cir[94] <=32'h3F7FE00D;
	Vec_Kappa_Cir[95] <=32'h3F7FE78B;
	Vec_Kappa_Cir[96] <=32'h3F7FFAE9;
	Vec_Kappa_Cir[97] <=32'h3F7FFC7A;
	Vec_Kappa_Cir[98] <=32'h3F7FFD6B;
	Vec_Kappa_Cir[99] <=32'h3F7FFE08;
	Vec_Kappa_Cir[100] <=32'h3F7FF808;
	Vec_Kappa_Cir[101] <=32'h3F7FFA7A;
	Vec_Kappa_Cir[102] <=32'h3F7FFBF3;
	Vec_Kappa_Cir[103] <=32'h3F7FFCE8;
	Vec_Kappa_Cir[104] <=32'h3F7FF483;
	Vec_Kappa_Cir[105] <=32'h3F7FF808;
	Vec_Kappa_Cir[106] <=32'h3F7FFA27;
	Vec_Kappa_Cir[107] <=32'h3F7FFB88;
	Vec_Kappa_Cir[108] <=32'h3F7FF05B;
	Vec_Kappa_Cir[109] <=32'h3F7FF525;
	Vec_Kappa_Cir[110] <=32'h3F7FF808;
	Vec_Kappa_Cir[111] <=32'h3F7FF9E8;
	Vec_Kappa_Cir[112] <=32'h3F7FFEC0;
	Vec_Kappa_Cir[113] <=32'h3F7FFF24;
	Vec_Kappa_Cir[114] <=32'h3F7FFF61;
	Vec_Kappa_Cir[115] <=32'h3F7FFF88;
	Vec_Kappa_Cir[116] <=32'h3F7FFE08;
	Vec_Kappa_Cir[117] <=32'h3F7FFEA4;
	Vec_Kappa_Cir[118] <=32'h3F7FFF03;
	Vec_Kappa_Cir[119] <=32'h3F7FFF40;
	Vec_Kappa_Cir[120] <=32'h3F7FFD26;
	Vec_Kappa_Cir[121] <=32'h3F7FFE08;
	Vec_Kappa_Cir[122] <=32'h3F7FFE90;
	Vec_Kappa_Cir[123] <=32'h3F7FFEE8;
	Vec_Kappa_Cir[124] <=32'h3F7FFC1C;
	Vec_Kappa_Cir[125] <=32'h3F7FFD4F;
	Vec_Kappa_Cir[126] <=32'h3F7FFE08;
	Vec_Kappa_Cir[127] <=32'h3F7FFE80;
	Vec_Kappa_Cir[128] <=32'h3F7FFFB6;
	Vec_Kappa_Cir[129] <=32'h3F7FFFCF;
	Vec_Kappa_Cir[130] <=32'h3F7FFFDE;
	Vec_Kappa_Cir[131] <=32'h3F7FFFE8;
	Vec_Kappa_Cir[132] <=32'h3F7FFF88;
	Vec_Kappa_Cir[133] <=32'h3F7FFFAF;
	Vec_Kappa_Cir[134] <=32'h3F7FFFC7;
	Vec_Kappa_Cir[135] <=32'h3F7FFFD6;
	Vec_Kappa_Cir[136] <=32'h3F7FFF4F;
	Vec_Kappa_Cir[137] <=32'h3F7FFF88;
	Vec_Kappa_Cir[138] <=32'h3F7FFFAA;
	Vec_Kappa_Cir[139] <=32'h3F7FFFC0;
	Vec_Kappa_Cir[140] <=32'h3F7FFF0D;
	Vec_Kappa_Cir[141] <=32'h3F7FFF5A;
	Vec_Kappa_Cir[142] <=32'h3F7FFF88;
	Vec_Kappa_Cir[143] <=32'h3F7FFFA6;
	Vec_Kappa_Cir[144] <=32'h3F7FFFF3;
	Vec_Kappa_Cir[145] <=32'h3F7FFFFA;
	Vec_Kappa_Cir[146] <=32'h3F7FFFFD;
	Vec_Kappa_Cir[147] <=32'h3F800000;
	Vec_Kappa_Cir[148] <=32'h3F7FFFE8;
	Vec_Kappa_Cir[149] <=32'h3F7FFFF2;
	Vec_Kappa_Cir[150] <=32'h3F7FFFF8;
	Vec_Kappa_Cir[151] <=32'h3F7FFFFB;
	Vec_Kappa_Cir[152] <=32'h3F7FFFDA;
	Vec_Kappa_Cir[153] <=32'h3F7FFFE8;
	Vec_Kappa_Cir[154] <=32'h3F7FFFF0;
	Vec_Kappa_Cir[155] <=32'h3F7FFFF6;
	Vec_Kappa_Cir[156] <=32'h3F7FFFC9;
	Vec_Kappa_Cir[157] <=32'h3F7FFFDC;
	Vec_Kappa_Cir[158] <=32'h3F7FFFE8;
	Vec_Kappa_Cir[159] <=32'h3F7FFFEF;
	Vec_Kappa_Cir[160] <=32'h3F800001;
	Vec_Kappa_Cir[161] <=32'h3F800002;
	Vec_Kappa_Cir[162] <=32'h3F800002;
	Vec_Kappa_Cir[163] <=32'h3F800003;
	Vec_Kappa_Cir[164] <=32'h3F800000;
	Vec_Kappa_Cir[165] <=32'h3F800001;
	Vec_Kappa_Cir[166] <=32'h3F800002;
	Vec_Kappa_Cir[167] <=32'h3F800002;
	Vec_Kappa_Cir[168] <=32'h3F7FFFFC;
	Vec_Kappa_Cir[169] <=32'h3F800000;
	Vec_Kappa_Cir[170] <=32'h3F800001;
	Vec_Kappa_Cir[171] <=32'h3F800001;
	Vec_Kappa_Cir[172] <=32'h3F7FFFF8;
	Vec_Kappa_Cir[173] <=32'h3F7FFFFD;
	Vec_Kappa_Cir[174] <=32'h3F800000;
	Vec_Kappa_Cir[175] <=32'h3F800001;
	Vec_Kappa_Cir[176] <=32'h3F800003;
	Vec_Kappa_Cir[177] <=32'h3F800003;
	Vec_Kappa_Cir[178] <=32'h3F800003;
	Vec_Kappa_Cir[179] <=32'h3F800003;
	Vec_Kappa_Cir[180] <=32'h3F800003;
	Vec_Kappa_Cir[181] <=32'h3F800003;
	Vec_Kappa_Cir[182] <=32'h3F800003;
	Vec_Kappa_Cir[183] <=32'h3F800003;
	Vec_Kappa_Cir[184] <=32'h3F800002;
	Vec_Kappa_Cir[185] <=32'h3F800003;
	Vec_Kappa_Cir[186] <=32'h3F800003;
	Vec_Kappa_Cir[187] <=32'h3F800003;
	Vec_Kappa_Cir[188] <=32'h3F800002;
	Vec_Kappa_Cir[189] <=32'h3F800002;
	Vec_Kappa_Cir[190] <=32'h3F800003;
	Vec_Kappa_Cir[191] <=32'h3F800003;
	Vec_Kappa_Cir[192] <=32'h3F800004;
	Vec_Kappa_Cir[193] <=32'h3F800004;
	Vec_Kappa_Cir[194] <=32'h3F800004;
	Vec_Kappa_Cir[195] <=32'h3F800004;
	Vec_Kappa_Cir[196] <=32'h3F800003;
	Vec_Kappa_Cir[197] <=32'h3F800004;
	Vec_Kappa_Cir[198] <=32'h3F800004;
	Vec_Kappa_Cir[199] <=32'h3F800004;
	Vec_Kappa_Cir[200] <=32'h3F800003;
	Vec_Kappa_Cir[201] <=32'h3F800003;
	Vec_Kappa_Cir[202] <=32'h3F800004;
	Vec_Kappa_Cir[203] <=32'h3F800004;
	Vec_Kappa_Cir[204] <=32'h3F800003;
	Vec_Kappa_Cir[205] <=32'h3F800003;
	Vec_Kappa_Cir[206] <=32'h3F800003;
	Vec_Kappa_Cir[207] <=32'h3F800004;
	Vec_Kappa_Cir[208] <=32'h3F800004;
	Vec_Kappa_Cir[209] <=32'h3F800004;
	Vec_Kappa_Cir[210] <=32'h3F800004;
	Vec_Kappa_Cir[211] <=32'h3F800004;
	Vec_Kappa_Cir[212] <=32'h3F800004;
	Vec_Kappa_Cir[213] <=32'h3F800004;
	Vec_Kappa_Cir[214] <=32'h3F800004;
	Vec_Kappa_Cir[215] <=32'h3F800004;
	Vec_Kappa_Cir[216] <=32'h3F800004;
	Vec_Kappa_Cir[217] <=32'h3F800004;
	Vec_Kappa_Cir[218] <=32'h3F800004;
	Vec_Kappa_Cir[219] <=32'h3F800004;
	Vec_Kappa_Cir[220] <=32'h3F800004;
	Vec_Kappa_Cir[221] <=32'h3F800004;
	Vec_Kappa_Cir[222] <=32'h3F800004;
	Vec_Kappa_Cir[223] <=32'h3F800004;
	Vec_Kappa_Cir[224] <=32'h3F800004;
	Vec_Kappa_Cir[225] <=32'h3F800004;
	Vec_Kappa_Cir[226] <=32'h3F800004;
	Vec_Kappa_Cir[227] <=32'h3F800004;
	Vec_Kappa_Cir[228] <=32'h3F800004;
	Vec_Kappa_Cir[229] <=32'h3F800004;
	Vec_Kappa_Cir[230] <=32'h3F800004;
	Vec_Kappa_Cir[231] <=32'h3F800004;
	Vec_Kappa_Cir[232] <=32'h3F800004;
	Vec_Kappa_Cir[233] <=32'h3F800004;
	Vec_Kappa_Cir[234] <=32'h3F800004;
	Vec_Kappa_Cir[235] <=32'h3F800004;
	Vec_Kappa_Cir[236] <=32'h3F800004;
	Vec_Kappa_Cir[237] <=32'h3F800004;
	Vec_Kappa_Cir[238] <=32'h3F800004;
	Vec_Kappa_Cir[239] <=32'h3F800004;
	Vec_Kappa_Cir[240] <=32'h3F800004;
	Vec_Kappa_Cir[241] <=32'h3F800004;
	Vec_Kappa_Cir[242] <=32'h3F800004;
	Vec_Kappa_Cir[243] <=32'h3F800004;
	Vec_Kappa_Cir[244] <=32'h3F800004;
	Vec_Kappa_Cir[245] <=32'h3F800004;
	Vec_Kappa_Cir[246] <=32'h3F800004;
	Vec_Kappa_Cir[247] <=32'h3F800004;
	Vec_Kappa_Cir[248] <=32'h3F800004;
	Vec_Kappa_Cir[249] <=32'h3F800004;
	Vec_Kappa_Cir[250] <=32'h3F800004;
	Vec_Kappa_Cir[251] <=32'h3F800004;
	Vec_Kappa_Cir[252] <=32'h3F800004;
	Vec_Kappa_Cir[253] <=32'h3F800004;
	Vec_Kappa_Cir[254] <=32'h3F800004;
	Vec_Kappa_Cir[255] <=32'h3F800004;
	
	//Linear vectoring delta
	LinVec_Delta[0] <=32'h3F70F10B;
	LinVec_Delta[1] <=32'h3F638E53;
	LinVec_Delta[2] <=32'h3F579450;
	LinVec_Delta[3] <=32'h3F4CCCE7;
	LinVec_Delta[4] <=32'h3F430C4B;
	LinVec_Delta[5] <=32'h3F3A2EA5;
	LinVec_Delta[6] <=32'h3F32165C;
	LinVec_Delta[7] <=32'h3F2AAAC4;
	LinVec_Delta[8] <=32'h3F23D724;
	LinVec_Delta[9] <=32'h3F1D89F2;
	LinVec_Delta[10] <=32'h3F17B43F;
	LinVec_Delta[11] <=32'h3F12493E;
	LinVec_Delta[12] <=32'h3F0D3DE4;
	LinVec_Delta[13] <=32'h3F0888A2;
	LinVec_Delta[14] <=32'h3F042121;
	LinVec_Delta[15] <=32'h3F000019;
	LinVec_Delta[16] <=32'h3F80000D;
	LinVec_Delta[17] <=32'h3F71C737;
	LinVec_Delta[18] <=32'h3F650D93;
	LinVec_Delta[19] <=32'h3F5999B4;
	LinVec_Delta[20] <=32'h3F4F3D0E;
	LinVec_Delta[21] <=32'h3F45D18E;
	LinVec_Delta[22] <=32'h3F3D37C1;
	LinVec_Delta[23] <=32'h3F35556F;
	LinVec_Delta[24] <=32'h3F2E1494;
	LinVec_Delta[25] <=32'h3F276290;
	LinVec_Delta[26] <=32'h3F212F82;
	LinVec_Delta[27] <=32'h3F1B6DD0;
	LinVec_Delta[28] <=32'h3F1611C1;
	LinVec_Delta[29] <=32'h3F11112A;
	LinVec_Delta[30] <=32'h3F0C6332;
	LinVec_Delta[31] <=32'h3F080019;
	LinVec_Delta[32] <=32'h3F878795;
	LinVec_Delta[33] <=32'h3F80000D;
	LinVec_Delta[34] <=32'h3F7286D7;
	LinVec_Delta[35] <=32'h3F666681;
	LinVec_Delta[36] <=32'h3F5B6DD1;
	LinVec_Delta[37] <=32'h3F517477;
	LinVec_Delta[38] <=32'h3F485925;
	LinVec_Delta[39] <=32'h3F40001A;
	LinVec_Delta[40] <=32'h3F385205;
	LinVec_Delta[41] <=32'h3F313B2D;
	LinVec_Delta[42] <=32'h3F2AAAC4;
	LinVec_Delta[43] <=32'h3F249263;
	LinVec_Delta[44] <=32'h3F1EE59E;
	LinVec_Delta[45] <=32'h3F1999B3;
	LinVec_Delta[46] <=32'h3F14A543;
	LinVec_Delta[47] <=32'h3F100019;
	LinVec_Delta[48] <=32'h3F8F0F1C;
	LinVec_Delta[49] <=32'h3F871C7F;
	LinVec_Delta[50] <=32'h3F80000D;
	LinVec_Delta[51] <=32'h3F73334D;
	LinVec_Delta[52] <=32'h3F679E94;
	LinVec_Delta[53] <=32'h3F5D1760;
	LinVec_Delta[54] <=32'h3F537A89;
	LinVec_Delta[55] <=32'h3F4AAAC4;
	LinVec_Delta[56] <=32'h3F428F76;
	LinVec_Delta[57] <=32'h3F3B13CB;
	LinVec_Delta[58] <=32'h3F342607;
	LinVec_Delta[59] <=32'h3F2DB6F5;
	LinVec_Delta[60] <=32'h3F27B97A;
	LinVec_Delta[61] <=32'h3F22223B;
	LinVec_Delta[62] <=32'h3F1CE753;
	LinVec_Delta[63] <=32'h3F180019;
	LinVec_Delta[64] <=32'h3F9696A4;
	LinVec_Delta[65] <=32'h3F8E38F1;
	LinVec_Delta[66] <=32'h3F86BCAF;
	LinVec_Delta[67] <=32'h3F80000D;
	LinVec_Delta[68] <=32'h3F73CF57;
	LinVec_Delta[69] <=32'h3F68BA49;
	LinVec_Delta[70] <=32'h3F5E9BED;
	LinVec_Delta[71] <=32'h3F55556F;
	LinVec_Delta[72] <=32'h3F4CCCE6;
	LinVec_Delta[73] <=32'h3F44EC68;
	LinVec_Delta[74] <=32'h3F3DA149;
	LinVec_Delta[75] <=32'h3F36DB87;
	LinVec_Delta[76] <=32'h3F308D57;
	LinVec_Delta[77] <=32'h3F2AAAC4;
	LinVec_Delta[78] <=32'h3F252964;
	LinVec_Delta[79] <=32'h3F200019;
	LinVec_Delta[80] <=32'h3F9E1E2B;
	LinVec_Delta[81] <=32'h3F955562;
	LinVec_Delta[82] <=32'h3F8D7950;
	LinVec_Delta[83] <=32'h3F866673;
	LinVec_Delta[84] <=32'h3F80000D;
	LinVec_Delta[85] <=32'h3F745D31;
	LinVec_Delta[86] <=32'h3F69BD52;
	LinVec_Delta[87] <=32'h3F60001A;
	LinVec_Delta[88] <=32'h3F570A57;
	LinVec_Delta[89] <=32'h3F4EC506;
	LinVec_Delta[90] <=32'h3F471C8B;
	LinVec_Delta[91] <=32'h3F40001A;
	LinVec_Delta[92] <=32'h3F396134;
	LinVec_Delta[93] <=32'h3F33334D;
	LinVec_Delta[94] <=32'h3F2D6B74;
	LinVec_Delta[95] <=32'h3F280019;
	LinVec_Delta[96] <=32'h3FA5A5B3;
	LinVec_Delta[97] <=32'h3F9C71D4;
	LinVec_Delta[98] <=32'h3F9435F2;
	LinVec_Delta[99] <=32'h3F8CCCDA;
	LinVec_Delta[100] <=32'h3F86186E;
	LinVec_Delta[101] <=32'h3F80000D;
	LinVec_Delta[102] <=32'h3F74DEB6;
	LinVec_Delta[103] <=32'h3F6AAAC5;
	LinVec_Delta[104] <=32'h3F6147C8;
	LinVec_Delta[105] <=32'h3F589DA4;
	LinVec_Delta[106] <=32'h3F5097CE;
	LinVec_Delta[107] <=32'h3F4924AC;
	LinVec_Delta[108] <=32'h3F423511;
	LinVec_Delta[109] <=32'h3F3BBBD5;
	LinVec_Delta[110] <=32'h3F35AD85;
	LinVec_Delta[111] <=32'h3F300019;
	LinVec_Delta[112] <=32'h3FAD2D3B;
	LinVec_Delta[113] <=32'h3FA38E46;
	LinVec_Delta[114] <=32'h3F9AF294;
	LinVec_Delta[115] <=32'h3F933340;
	LinVec_Delta[116] <=32'h3F8C30D0;
	LinVec_Delta[117] <=32'h3F85D181;
	LinVec_Delta[118] <=32'h3F80000D;
	LinVec_Delta[119] <=32'h3F75556F;
	LinVec_Delta[120] <=32'h3F6B8539;
	LinVec_Delta[121] <=32'h3F627641;
	LinVec_Delta[122] <=32'h3F5A1310;
	LinVec_Delta[123] <=32'h3F52493E;
	LinVec_Delta[124] <=32'h3F4B08ED;
	LinVec_Delta[125] <=32'h3F44445E;
	LinVec_Delta[126] <=32'h3F3DEF95;
	LinVec_Delta[127] <=32'h3F380019;
	LinVec_Delta[128] <=32'h3FB4B4C2;
	LinVec_Delta[129] <=32'h3FAAAAB8;
	LinVec_Delta[130] <=32'h3FA1AF36;
	LinVec_Delta[131] <=32'h3F9999A7;
	LinVec_Delta[132] <=32'h3F924932;
	LinVec_Delta[133] <=32'h3F8BA2F6;
	LinVec_Delta[134] <=32'h3F8590BF;
	LinVec_Delta[135] <=32'h3F80000D;
	LinVec_Delta[136] <=32'h3F75C2A9;
	LinVec_Delta[137] <=32'h3F6C4EDF;
	LinVec_Delta[138] <=32'h3F638E53;
	LinVec_Delta[139] <=32'h3F5B6DD1;
	LinVec_Delta[140] <=32'h3F53DCCA;
	LinVec_Delta[141] <=32'h3F4CCCE6;
	LinVec_Delta[142] <=32'h3F4631A6;
	LinVec_Delta[143] <=32'h3F400019;
	LinVec_Delta[144] <=32'h3FBC3C4A;
	LinVec_Delta[145] <=32'h3FB1C72A;
	LinVec_Delta[146] <=32'h3FA86BD7;
	LinVec_Delta[147] <=32'h3FA0000D;
	LinVec_Delta[148] <=32'h3F986193;
	LinVec_Delta[149] <=32'h3F91746A;
	LinVec_Delta[150] <=32'h3F8B2171;
	LinVec_Delta[151] <=32'h3F855562;
	LinVec_Delta[152] <=32'h3F80000D;
	LinVec_Delta[153] <=32'h3F76277C;
	LinVec_Delta[154] <=32'h3F6D0995;
	LinVec_Delta[155] <=32'h3F649263;
	LinVec_Delta[156] <=32'h3F5CB0A7;
	LinVec_Delta[157] <=32'h3F55556F;
	LinVec_Delta[158] <=32'h3F4E73B6;
	LinVec_Delta[159] <=32'h3F480019;
	LinVec_Delta[160] <=32'h3FC3C3D1;
	LinVec_Delta[161] <=32'h3FB8E39C;
	LinVec_Delta[162] <=32'h3FAF2879;
	LinVec_Delta[163] <=32'h3FA66674;
	LinVec_Delta[164] <=32'h3F9E79F5;
	LinVec_Delta[165] <=32'h3F9745DE;
	LinVec_Delta[166] <=32'h3F90B223;
	LinVec_Delta[167] <=32'h3F8AAAB7;
	LinVec_Delta[168] <=32'h3F851EC5;
	LinVec_Delta[169] <=32'h3F80000D;
	LinVec_Delta[170] <=32'h3F7684D7;
	LinVec_Delta[171] <=32'h3F6DB6F5;
	LinVec_Delta[172] <=32'h3F658484;
	LinVec_Delta[173] <=32'h3F5DDDF7;
	LinVec_Delta[174] <=32'h3F56B5C7;
	LinVec_Delta[175] <=32'h3F500019;
	LinVec_Delta[176] <=32'h3FCB4B59;
	LinVec_Delta[177] <=32'h3FC0000D;
	LinVec_Delta[178] <=32'h3FB5E51B;
	LinVec_Delta[179] <=32'h3FACCCDA;
	LinVec_Delta[180] <=32'h3FA49256;
	LinVec_Delta[181] <=32'h3F9D1753;
	LinVec_Delta[182] <=32'h3F9642D5;
	LinVec_Delta[183] <=32'h3F90000D;
	LinVec_Delta[184] <=32'h3F8A3D7D;
	LinVec_Delta[185] <=32'h3F84EC5B;
	LinVec_Delta[186] <=32'h3F80000D;
	LinVec_Delta[187] <=32'h3F76DB87;
	LinVec_Delta[188] <=32'h3F6E5860;
	LinVec_Delta[189] <=32'h3F666680;
	LinVec_Delta[190] <=32'h3F5EF7D8;
	LinVec_Delta[191] <=32'h3F58001A;
	LinVec_Delta[192] <=32'h3FD2D2E0;
	LinVec_Delta[193] <=32'h3FC71C7F;
	LinVec_Delta[194] <=32'h3FBCA1BC;
	LinVec_Delta[195] <=32'h3FB33340;
	LinVec_Delta[196] <=32'h3FAAAAB8;
	LinVec_Delta[197] <=32'h3FA2E8C7;
	LinVec_Delta[198] <=32'h3F9BD387;
	LinVec_Delta[199] <=32'h3F955562;
	LinVec_Delta[200] <=32'h3F8F5C36;
	LinVec_Delta[201] <=32'h3F89D8AA;
	LinVec_Delta[202] <=32'h3F84BDAE;
	LinVec_Delta[203] <=32'h3F80000D;
	LinVec_Delta[204] <=32'h3F772C3D;
	LinVec_Delta[205] <=32'h3F6EEF09;
	LinVec_Delta[206] <=32'h3F6739E8;
	LinVec_Delta[207] <=32'h3F60001A;
	LinVec_Delta[208] <=32'h3FDA5A68;
	LinVec_Delta[209] <=32'h3FCE38F1;
	LinVec_Delta[210] <=32'h3FC35E5E;
	LinVec_Delta[211] <=32'h3FB999A7;
	LinVec_Delta[212] <=32'h3FB0C319;
	LinVec_Delta[213] <=32'h3FA8BA3C;
	LinVec_Delta[214] <=32'h3FA16439;
	LinVec_Delta[215] <=32'h3F9AAAB8;
	LinVec_Delta[216] <=32'h3F947AEE;
	LinVec_Delta[217] <=32'h3F8EC4F9;
	LinVec_Delta[218] <=32'h3F897B4F;
	LinVec_Delta[219] <=32'h3F849256;
	LinVec_Delta[220] <=32'h3F80000D;
	LinVec_Delta[221] <=32'h3F777791;
	LinVec_Delta[222] <=32'h3F6F7BF9;
	LinVec_Delta[223] <=32'h3F68001A;
	LinVec_Delta[224] <=32'h3FE1E1F0;
	LinVec_Delta[225] <=32'h3FD55563;
	LinVec_Delta[226] <=32'h3FCA1B00;
	LinVec_Delta[227] <=32'h3FC0000D;
	LinVec_Delta[228] <=32'h3FB6DB7B;
	LinVec_Delta[229] <=32'h3FAE8BB0;
	LinVec_Delta[230] <=32'h3FA6F4EC;
	LinVec_Delta[231] <=32'h3FA0000D;
	LinVec_Delta[232] <=32'h3F9999A6;
	LinVec_Delta[233] <=32'h3F93B148;
	LinVec_Delta[234] <=32'h3F8E38F0;
	LinVec_Delta[235] <=32'h3F89249F;
	LinVec_Delta[236] <=32'h3F8469FB;
	LinVec_Delta[237] <=32'h3F80000D;
	LinVec_Delta[238] <=32'h3F77BE09;
	LinVec_Delta[239] <=32'h3F70001A;
	LinVec_Delta[240] <=32'h3FE96977;
	LinVec_Delta[241] <=32'h3FDC71D5;
	LinVec_Delta[242] <=32'h3FD0D7A2;
	LinVec_Delta[243] <=32'h3FC66674;
	LinVec_Delta[244] <=32'h3FBCF3DC;
	LinVec_Delta[245] <=32'h3FB45D24;
	LinVec_Delta[246] <=32'h3FAC859E;
	LinVec_Delta[247] <=32'h3FA55562;
	LinVec_Delta[248] <=32'h3F9EB85F;
	LinVec_Delta[249] <=32'h3F989D97;
	LinVec_Delta[250] <=32'h3F92F692;
	LinVec_Delta[251] <=32'h3F8DB6E8;
	LinVec_Delta[252] <=32'h3F88D3E9;
	LinVec_Delta[253] <=32'h3F844451;
	LinVec_Delta[254] <=32'h3F80000D;
	LinVec_Delta[255] <=32'h3F78001A;

end

else begin
	
	x_FSM2 			<= x_FSM1;
	y_FSM2 			<= y_FSM1;
	z_FSM2 			<= z_FSM1;
	k_FSM2			<= k_FSM1;
	operation_FSM2 <= operation_FSM1;
	mode_FSM2		<= mode_FSM1;
	InsTagFSMOut  <= InsTagFSM1Out;
	NatLogFlagout_FSM <= NatLogFlagout_FSM1;
	
	case(state_FSM2)
	
	Circular_Rotation_with_table:
	begin
		if (enable_LUT == LUT_Rotation) begin
			theta_FSM2[31]   <= ~z_FSM1[31];
			delta_FSM2[31]   <= ~z_FSM1[31];
			theta_FSM2[30:0] <= Rot_Theta[address][30:0];
			delta_FSM2[30:0] <= Rot_Delta_Cir[address][30:0];
			kappa_FSM2 <= Rot_Kappa_Cir[address];
		end
	end
	
	Hyperbolic_Rotation_with_table:
	begin
		if (enable_LUT == LUT_Rotation) begin
			theta_FSM2[31]   <= ~z_FSM1[31];
			delta_FSM2[31]   <= ~z_FSM1[31];
			theta_FSM2[30:0] <= Rot_Theta[address][30:0];
			delta_FSM2[30:0] <= Rot_Delta_Hyper[address][30:0];
			kappa_FSM2 <= Rot_Kappa_Hyper[address];
		end
	end

	Linear_Vectoring:
	begin
		if (enable_LUT == LUT_LinVec) begin
			delta_FSM2[22:0]  <= LinVec_Delta[address][22:0];
			delta_FSM2[30:23] <= LinVec_Delta[address][30:23] + exponent;
			delta_FSM2[31] 	<= LinVec_Delta[address][31];
			theta_FSM2[22:0]  <= LinVec_Delta[address][22:0];
			theta_FSM2[30:23] <= LinVec_Delta[address][30:23] + exponent;
			theta_FSM2[31] 	<= LinVec_Delta[address][31];
			kappa_FSM2			<= 32'h3F800004;
		end
	end
	
	Vectoring_by_small_fraction:
	begin
		if (enable_LUT == LUT_LinVec) begin
			delta_FSM2[22:0]  <= LinVec_Delta[address][22:0];
			delta_FSM2[30:23] <= LinVec_Delta[address][30:23] + exponent;
			delta_FSM2[31] 	<= LinVec_Delta[address][31];
			theta_FSM2[22:0]  <= LinVec_Delta[address][22:0];
			theta_FSM2[30:23] <= LinVec_Delta[address][30:23] + exponent;
			theta_FSM2[31] 	<= LinVec_Delta[address][31];
			kappa_FSM2			<= 32'h3F800004;
		end		
	end
	
	Circular_Vectoring_with_table:
	begin
		if (enable_LUT == LUT_Vectoring)begin
			theta_FSM2 			<= Vec_Theta_Cir[address];
			delta_FSM2			<= Vec_Delta[address];
			kappa_FSM2			<= Vec_Kappa_Cir[address];
		end
	end
	
	Hyperbolic_Vectoring_with_table:
	begin
		if (enable_LUT == LUT_Vectoring)begin
			theta_FSM2 			<= Vec_Theta_Hyper[address];
			delta_FSM2			<= Vec_Delta[address];
			kappa_FSM2			<= Vec_Kappa_Hyper[address];
		end
	end
	
	Idle_state:
	begin
		kappa_FSM2 				<= kappa_FSM1;
		delta_FSM2				<= delta_FSM1;
		theta_FSM2				<= theta_FSM1;
	end
	
	endcase
end
end
endmodule
