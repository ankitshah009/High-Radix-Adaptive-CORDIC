`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date:    20:06:14 11/04/2014 
// Design Name: 
// Module Name:    HCORDIC-Main 
// Project Name: 
// Target Devices: 
// Tool versions: 
// Description: 
//
// Dependencies: 
//
// Revision: 
// Revision 0.01 - File Created
// Additional Comments: 
//
//////////////////////////////////////////////////////////////////////////////////
module HCORDIC-Main(
    input [31:0] x_input,
    input [31:0] y_input,
    input [31:0] z_input,
    input clock,
    input mode,
    input operation,
    output [31:0] x_out,
    output [31:0] y_out,
    output [31:0] z_out,
    input load,
    input next
    );


endmodule
